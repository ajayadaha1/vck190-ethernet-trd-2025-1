`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
VrNh7bjPAtWwAmHLdNvs7XEqkUnMigEXGK+tVeTQQ/TzQBessxFdhp1tw+y7ozn8RcYW77GnU2W1
Visba6TKbjgZtujb4C/JQmdjNbzRPvdE27Av27pJEKMToJFORfFT+zPLEOoyhNIdx3Js6rqZ3f2b
54gXm3i+6LFZowSh/7Pag9mb3rT4wEZPNWwHaM4PVGXcAH/rmDNxpB0+baxk8vM/jnOptKyyEvco
+KpDhR22m6rUvOCE02LxIe8uX3tK32pwNaGCBcuEfeaHjM/OFfnh0UiFAE2EpgQcRIWwTiOcpTN/
cexCsDFURa7SBn9SpwPsc6WUgDtJ6bw+2/rLBw==
`pragma protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
uTesPuubgqWhsNh2+VhVeZ6O2WO19nLo/T1Kxcp3MWhPCucfKCcTibOypmCt4Lww+8WBBVwaYbg5
ULDumjjdu+uxXX7Yyex0C2OlbklEc6WSdyrbX8k6BQkO81PdWQ3N/Tvfzgds4Cyun5a/gdwVgJ13
HB77u0lWpo2pT0UadhECvERsD2bntp/0nT+C4uzv+CvcYMt4Fr87zOe+DoEBz8FzWk9+561yR/kR
xxRDdl20DZ8rRvglcIDsYRMuX6HALrunIZQK4WKiS1Ub5TUiNbI1uVeda/MJ4QDEhc/Y0GBCPSi/
RdrUAlzUIu/7XK8H3QgcwjChGteNAkK53ckUpA==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
RlUHmAm5AwnStJEa04JA0lAjR2wMpFoE8RNr/1FxXIj6zizuNPFpAJhDZre0nFlLZPUjuImgXv+0
LNclH64nSA==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
XFo5EAaxKwGtCu5vmN8gUas4DMRa+pHlK4cDVBF18JRNwbtJIrjbCZAtp+AMF+gUjAJ/5oJstlMA
EMPhtZrx38jfOUU2Mmywb6ZvIvI+dkg4M5vtQjt1XLN0O8nzZc/hWSyk9a2ZgVZX0c7L5rcGku7L
zQhR/4NhO3yKQarP7oQ93FvrBm5XYo/Za3Nzm17vJEOqsJ7pePAoq3F2wBElBkAG8WSwsmcfmio3
3wmheKxVbEVeQUyIUZywjJ3td2MnBnxy8/gTwTvB2eONp7hR1W04Ggj7BeG3HOGKkTwEe3pCWXRl
bYZtc56FvUitGhhlXjbRP8Q5o9M2j0bqlQKIkQ==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
K9FRPo7Ddj9rzV0Zd9kHO2Vd5Y8VgRBTQ8whDExoCydRri315aEcPRmgM1QzOV7EQhxAMw29TOPS
I85qhYEFRffVrweT5FRRNjPyNLIlBeHo7CFTbpBZeSMDqIz0yZ4uErMqgTNofANDb3q3xxkzE5w0
N/w0O7ffhcQ7Z/iyY7I=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OuJn0UR3AQAvVKWKq/HzCJMB3u21GVREGgBioYtpxg8I6oWeCg9IO8dBndQo2P8y7laXQ+WYh7z9
JeealXbtwSJLn3L3RvjHtA1rT0Y03LoWC2P/3vYsmXvFZQvVYM43+SzTVhhwEfDUJ6y6nh8QVso7
nCUUp0Ewx8OKvjAqbJBmBQ0jpTYFN9/WS4ZZuUG/IH95URH5i/o5hFFGvHD8MYuKfIZNKo+3H691
tt62kzCr0diVOjMBlN8NFN/YL7ID8rzSQ93Se655lL2nk73yUlvdN+mIqPbu0GXbqAwFWqZnDzgL
YqIoVfuB5ISq5QXMAWsoMpN21Ugzrs2v98ryvQ==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
t0Y4+mUnuvt4CMcmeOMXyK+/kj7A1Yf6NW/x2nEZIwOyLU90qMUCloC1DSZaCXX/xpbzz1PlO7oJ
nTzqlMLhMb83BDBkeHvX+BTCU4se8NoI2GKlCvysW/CLvom9uuPE9Tn0QTbv1urzKVoVl/EiatZC
oWg1JDftrwfydzaL3OwEG/PeGs889kym2/UOyj1Fbn6aMwA44o788tnC8QSmNp3mIUNrmZZ+IqOx
wJcnG/VgZanUgRodmyIfaNmZZi8yqnVUduoOHC/JZgVQMQs9Q4wW3+GxpkGgrJzVqz7tSUDj7keT
z5KPPdi2D0qovwui8H0W1Y/b5UAQ5ryqDinPJg==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
uB+IfF7V/HDqA7+3E15U2WjuR9aNtr2gzwkShm7yKE+8sHg6il6bnMNJeLO0NyPnTIosyTMYaNZR
WzSJGhvh3HpgD5woUWE7gVAomxjoKbtDUgLu/VQTD3RCjkQg+Uddg3s8w+PZnPkj6CfP/mS9qaSb
XooNWdEl20W+zzt6srk=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nWMQTBfWtdFpCZ0CWPX4++z/5eraGLaln99q8Hoe5XCCVqtBzAgU3UKzRlZ290VSR5FHoF+VAZZU
ZvBPazGTPzXKFaJ7WN++iBm8y2lQ6W5LOhSOjjs0Psc7fET2wdHLO1EGWtjhy7kBZABXnvbhCJTJ
47W5m+h7ikJgTNwaLsl9U3uc8h51KsxDSRcSAksaC6pjw0yJGLCcytAzhwHM3mkeWuYaxUoe7ZoK
yGvwdtT6kyGiL38tD/4JBVCgUUzTJJ8UxNO+lBA4Khn4ejo+p8EQR54YIMZfRm38LjcGF81eG1PM
xD8wKeXhR3Z/tHcch51jMkmWrsxbtr+f1cWvlQ==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12800)
`pragma protect data_block
OEJgQdUiYYt+N0r7zKCecfkVMfAfOGUDO5yJC5jssBPXW0Zk3JDjWrF1etDjUIg77nvqVSZwF6Fn
vOvYfSqm4III+bYE1Ev/djD24fjBwwYWCQ7Ha2WtTFFcbvRlIjZElLkNZglXPlWm3+ukY5s4XJyC
CfBuYwprAPExnu9W2kkWpeUwApOih/+xMtKaDvJ1mVUr+WL1nEIMeSyPxADjpY1DVXWNPgggZjse
jRlvy3+ID6fpd1sLj2FJIfCN11QAcMgs2vkKkxeVHSX0j4k56EoXk8v0xg5dxeQHWsOfG82Jl1pE
QAGhDSMbln5s8FqER5d6tZGiEV/j/LByodLds+q32KtxDleDnV9meLMRgLVjhdOADwfyJ/pkQydU
ITwEP7BI6bNrJ9Q53Dxk3WwRX7yJXXgGPRNoiEd4c0I0/1SO7QMYrbqQ/U+wBLFS9ywPr0DZArMU
ITQLMicwEVACYPPAaUC+w9GpUUdSEg82TPF0laMsCA6OCXfW5S7RgVgb6VM5W4BUNe83VZqW4+t1
feNVSSfcSCXTlHbVpp2IOkW9Il/NZeRXH/aURCWubbSfq+ILSGWXdu9vIuCnXVSAOBkLTgQRjGu5
j8XFS8h1sjAdgFa6X4CHVItocWxgJEuVudilrZfU4o5DjtN5wo6p4pK5PWbV/pXyIVl1057vYKAR
A2FfgxxKtWZwr/65OaE404+hbGyYpCzFVKWZqPzb0pi7CGEN37xWOlXBR1raL8CtvAys5XOT7NPR
nRRQeK6QKWVMmZPNrnhiIgkYPDtpMmN+arSV4sxdZ6VG7ywiwMx6DLV4yLL56pjYAi72QqnTrrpC
jpiM+I1yKqyyTr6loASnjuzk5+wv1OfT6BezxhSxXwqrcymP1MXFHu5g5NOIZwgGo2fGe+DWQwdP
sKHHf/BGdkHIuiXkHsrsF6gfL8mp/mx4fqYIF1zre5tQq3EK3Z5cqrpj73rcLOQaYZXIj4EaF38T
4l4rUq8l3WQof1NUZyfvjnlTws1oVKd/KVtsxoAye8sWsWqsy10tnO0xbqU/yM8KvCfPTGtSIaSi
FpoZ39ICCsDzouFxLUqbni24aGlh+lo+kb7NJG2amAiUJHOWFT36/8Ag5VLeHhrn4l6ZkvllW/vV
h7USQVa0FMEU2B3mmrrm4QiDah1zixQVAHscU2BtM2JY+XlyvcSQObc/G1I44fcx4lOS55yhzmvB
+3D/4m+40A7Q6NN3kSfgZ8UIE+NGwCrpGkvj9mnEk9vCrnT1AjaO0vFum8UTUKQQsxFIx9s8CXFH
cZzZplM64tzd9XKv7/u13dlBfaySWvgrAIKrkNWIVVgj3VLelW9U0oPfGdB+CeQe4QStYW6guNX3
DkSz2xgFODHckniYO9Fx81ukTybAfvAGUHwt9sKMjKawPe6qMOawz+Z6rv1cYcuulFOHcnvxl6sq
za9ugYArhTO6IRMDYJo4fB1FSQBt7pNZFKet8HIGjicNncCt9l37c7rKk/xyfL1XSWWh3QcFCBa2
/a/uemtcpSK0WmgcF6o0DYDe0RztsAK/gOiBEZgcMK/pGJ12BTYEQpJEDXcMpCAFXt6jovoVLdCi
aPCaz9M4BDRZaLWzllWLn1k3pX4fF8wujSXBfDtkpKeLkKtdLFif379sMo34RvXd8Fnw06LrZe4W
1tTissAf78h0ZACICHAYxN1VI65eIAuj5aI+rIEFZuyIdtAnQWr9E9Sqi7Oc8tQFd1gVV97ltbGj
OMTEjUEnk+yb0lcPIzly7F4V9KW6dL+vTTvm+gQRBr+mRxhctWcMK+vAlk5emoNjiWv1ye6fQpL+
ilGFqCVXsFPMYilCnQ14Pe/t47Bf1NsMmXwjRXlou67FvOVpR8JkyuIoYcTl1v+Kun6f1U6AvjB7
/QOqdPEZHdEwe2VI7xZN+hFDnwny6uLuc+cxqn7BWEy4B33MRYbvDJ2iEy4KIMmqttTANyrzldwt
Qp1TgAPqrIjKCfanKRnBiWscanZ6gVggQUyFxt+06IheaQ0+5fUvbUA3zL3MZWYvEDCneQM4dpWi
yPRhKBWgQ/C8+soZXdZi/DLYUQVRM8wUvjVgX9UJVhyUoIPaY05wkdYyywLjGZJN12Vo/AEuK5vO
DJsPWAZPfqgeJHgiShOkkex1qZi34CCjBCMcu1PCewjWv/1mvbqNbqxKn7wl8gjkr12qhPsI7n+t
FfVJKxNtKoWGAoMbn/MzuW/Fsq3oWPmwFo2RVNqwceLDWU7MrA2OJpF9N0UAIt/KM0BpzW3NELzi
gXEDl3vGpG+eWJV1/MfvlduraU6zvzVR9D79arzDIe5tKJZgMQX6a7Wq84AI5/JPu7VOwzsAUyi5
nAuMAVtHD7LcIsbcfLAMeSnFE0O/Y8Ay1N09jwOa/cv/8C3P8naSojDlfq4UL20nhkN9hNdT/8J5
m+Hl8g4Lztmlyadr6WydNF4mRe20TLf/OeA9G5GLba50yunv8yvpUcM0u0nDDTXFdNs52LKAyh7I
QPnuP9GuWbXr5FeJ5lAsORpU5PuPRdZWoyfxDevBLo8z+43tMhgrXqn0ldBDSld61vMIR6Ojs/cH
Kzt1gvVMmH/K4s7+ecYCeuXm1ostYGf0vNllT+2DPfYn0ghBViDUxR8eP4ikGBzA+vO8EBn3WkZe
pClyrrVZsCgVUEkqWl5VZxokoVL7BI0IX9PmoD7uqpcaUc1lf+8oAyJ865pyHshxy4ZeZzDO/+1a
ILsQi8DUum8WYgHTqJm1Q12hGnlIGuTGq9E3ityrMOn5A0Ch1YWZgyhD+PezDOesz0RAh5K7l/6I
yH436VVtUIqi4zzyeO0Qm0ZrnEysSCsvj2MKWNPbaSzmI5i3hYcvJF2nQxwN2RrNzKrZD8aUY4od
iflOQcqbdLslUj60pYpDbE7aEdiAvQMwgm14EQnJkQgYWLi/IDgb5EwbitsTcYMGRe1yHVxCQ34v
D6a2L28FQJqySUMsVdeB5ONUkoOrcdY23gJfEWxQVRqr2ffdM+dwPvY1cvdXI7ZYV5kK+wp0u22Y
Q9VkGFyTDBoWiBZ0wwxMDctKASL1vs+CGRcCu4s4+gLxeewC+OGH6vqXZwK1fX8S57BKeBgv3I+k
NGjKA8legsj6SQ2uV6T3dfusZcmSFTlW9LTY6zgaUCnnSy+V6Bz0aOHXV0IpFExX78CTN8Ow5mjx
Qh2GmbvGOY1qUy9HdzoUekatM7YVC/nlwJ0i/ReDG6GX46X/ADFCPlehlbQCOpk5+TVvnM20DXSH
+GZGwKi9IAodCueQKQ5SZ950rVQMDUXlH46JAosUpboMc725WbUt6SLHWuLQLhudLaKvW+jJPBX/
O0s/7P2K1pQ3rHryB77KjMCWnRwr7Pj1DT5HuSG2YfxClKfS7OXDAvnUTqA58g4t3C0iMU5xw2PG
sQseq2vnve3FiuXT1H1hqANhX4Mp/zaoC1+vahDGyuk4LpqJlxf0uB2q2bnF/1gD+BN2us/VvhfZ
r/+Nie+eqGv8dpMRJNYLYMPLcnSlogMLU7XUX5O9lvPvwf1hn01t5lcX9Aclx1rZ4kGrejb4w4gF
xFnqjno5IzRxe/h6l33wIUqmEeU+2YydKjxekpU8dwPZDMjthb4xPoYvGHQmC0enwNkjCMHR1fIS
Vl8Es95LnO1ReC2a2nsdhLqbnUnzBlLyg29tUWtVcsnPLxLFSM0w69MZ/QF9lJhFCOop7RG1e87B
uYqJH6o+wuL8RwJan3fwXW1nkDdVvJ+d6lVJAOkMO+hzBLqg/SoCltzq69qzdH8tuI4DVOBGZPMv
Gcfmf7MFbFYMT6pRJdWxjqUniZVuaLN/pBwJ9ShG4Nxz83D8SY5vWfiqj7ZbjFw8sj5jfQrNRA6r
WhBmU1w/sgn4boK5EoaPfOCcxr2JSEQQXJfFv++2VC3EQyrcVnGa1mZ+e+rmDQM8jCU2dSpyp6Pd
R8ZqOUzYzsbjlr6Jt0lg3VO2To21DCI6uhIU8+/FMMQdpofyvygfKcr2Ax0hlO/1sykTB8vucB24
dcc+GArV+oDmJRq0BYpl/tWUkA5BDrr9IuwT82HjaeBKcPH8WB6onX2n9Ot8M5iTSbsx0JUYticj
N79CivsWuKDFom5IqeDmB78B6J+uekVvR272e8bU23dvoRXvnM2CcY+SKYTCnEFRtvjJB6tJAr4Z
3b0q2CIvGVuE/poIz/BX6J0M9qvLcupLUvzaywbYbIjGMHKIrNuqTctYjhAbvGEsFmkazAdSoeQj
SUx+3oI1f7PEFWEiRr+wUCb5JjVF++IjI7wfumb9xcQT4qYMldeNnSNTIteC7g/5Ftb3090pLOXF
BZ13US4/kFAcCPgUn35LKhga7aJTtoSD2xm5DtqugMAWSktYVvVo5fZhJEkzlbbbo739R3oiwuxB
6/UUX04U8I4S4X9UOIuhIabyqPbHTiLXH9dydehSsq15o4Ybu72Ov9MqVEL5ldnNZYU2LfJ4TDFB
7FUc3BWYkWa70VFd4KTOyZ4Ai1G+hX1VtF3kksQdN2cwlfHMI9uweLwxxsIVwJ1NC2t1cufcAq4j
1s/7yOv8lP+IXmd7YmBpB0UV1SHgnpGj6bWpAMqlA+qWEyTcJGXIhPPsD9/Mq9YsC/79rgiPBLlJ
IAy/qYI27BlCMZ14KQhddHnMBgdVvq2W/9F9ac33EB5wOvdYgAyc7eYKf7/iwfIa7XKPRmu2OypO
WG5rZE+VCyXlwhRRu5DAFTgxGfwvM8uwUh25JTsFrAqt87ZJihA91tnr6+j+P/fLieHNy77nyU8P
o00qqwlEA76mXCsXqd+YhvLA+QLN4nQKOkCdTL2rDW40hlxAep+G2mjzO3xe+xIw8O4Tv/bxNEfR
5j/0ZuR6aNHPuXS2b6sYcDaXvFX8fCsecwN9OoVMsEQX818vtFPcX4+CYLhNeVFNDOFrPXEtuWWy
g1c1dtA04EmJf6Ze7tPckgMsZm/v8IFRNPwUXIqMbMAmRLM7S9HF6W/t/RYLJE3tzhc2VCPUfZl7
EgQFsk5gvH0TciNgAGKGFJedqysPdjxlpYVxByZDGg1edQYlvrtlBYUJGPF0T6ua2eSy+1Jix1b6
yoeTMMRjQMQ5qYwWINeokHZ+MYPLeX+xN0B2UettM90TQsgqsG+PQ1rOjVFxC68Va2r0l0f0MYPd
Q5F4ViGCAe9Kddd6S/jgFcC6nbGvoRNkwNLe9FpkIz0Bvd42+senqJERsFmO8CPjb6ZUIqqJN+uU
enxLt/zQIEUu87E751o+ZAhh0y8xu2a5VuRwGCPt6JdUCF8NQaJdMTkA6ZfI1vARmqunMgEsCYHK
kefw3KBrGDjxd+huUgcQltZvJh9FNWU7eIIqnXDCqGrdI0sfissplhe31Lr4eqhGUM4DI7r0NLx6
fjwGd28V06wF4pkaPF3epyxpysrbvTTWX4J9FUtmTQDaP0ZEGvmcHpqiv0NGwtH508GZMuaqxlsV
pXYpUNbch2vDYmTdhifD95lc89U4Q1qkaagIRt5h5uYCVzXOm9g/QnwqZFefdKgqH9t3sf2D/JM0
unB9fqHdoLFKWvgY/Qz1NS6eI5uaBXb3nmi+JeEDHWV0on9eD7484d36bSnAAd5bjboeWZWFeg8r
Nx/JYBCuU4DSFYOyLVI9FNw0SUV5rb+d8RZRmleeKJkC2wuoHQlT/WekK4B+RrTcNtvaXf3BtPhc
D2TMEDRohgAF/SwCwWRtj1AqcAko8HSaOIqOewwkC8YaSwJWsUUqKtWY50jgIUBUEUAljZxjd7k4
so0Oa8Ntc9Mqf/K/29I1KJQTd9w7BUMso15pq/BijiVgf7mUgkYsEHHsqlVBAKi3zF7LxBYbJJop
WQj/+x5i0eZ6wq77Nk3xoR4TWkyq4BnLAdrbeJEvT2xBmuuVZFLxyLYu6l2Ymrb0U3RsQvvwhKSf
xYUYB56LzgzSddq0kU3Y7aXshl6lKAA8W8KgRoSz7iRKsuPbj6ESivviIsy4E0ziUChssEJJr4uc
9WQkbRCv1zXyhmujhX1Ei4Bso8rPf45ckq22/h6+7YVwpBcU3NFDF5q/YNlMYCbeKMEo3TNgAN0M
bTD7SSHzDpvjYCZaHghk3s0/NkNs+7BBjjIU1tJL5kEcNemfiVywfBXaewcxyEO1gRsNrVYvtEr8
wkcYncTd/5nKMONNDqGV8e2trUlzf+b/S6WM+rekjKQLKCQgUwjZHC76gvnpItHl5or86dRHeaaA
qjiKJVKT8jWX1HrYL67vsNZ9NMgy/OXUNNsfISYdn705Nb8GuXP0o6715jhzm42Nm7GL2+eZmt1R
5OOWV/xJuxEbWknPlLQeTpXd2aGFdt0hkaxhc5DyGYeeNjcTjeRDOrE+5ioc6mpal42uLAuJiARB
htd/rAf+zJeRpiO8xYb0R5EYKqAVS8NXW9upqRuuhR46lhOs1WUHrWZpQ3w6XFBfzlWpmk41lR3S
67auhY6JjrmMD+kGTbJCPGWIAvQFzqnVOkGZeZ8Nib/h+9iVS5JB/mtK77Ak0iY41QNpGQaNJBoT
Q/eYQ7rLpoZfSloA6HFgbqklHpAzo0l7ENe7gWgOKhcJBfmeylv2x3+LWit9lGNPystcwgCVLF9G
0ejlEq8ViuoMei+6/PLauFho1uhPMCkA0Qi4igl0oc8NW5yPz2TqABXYPmayX1XZJrAfLdPCRZJ0
t6FqR6p7VORcxEfbhkp6v3u2dFzJUh+idADPBlwKp8+C3H5cCc2i78iG3L3UhhvCuO64pVR9sBpc
MFw635pTGPODruI+1OKJC+zztbWNTrJpxK3vV1hX0FhLn4lLbuXLZ0ybvKJ6QiA/uEMJ/0orqNMu
yCgfxzDGOwSm34tIE3K9ZNfkS8YK3VBp3MClpTPP8yAeaCYsiL2XJ4CZOTFTKzA/WF1ugxcAuyGD
klRQTLtq6O5fEDTsrkPascnGgbE3+xLOfovcLRfffJ7n7gF0XYNVrS108TzrkZmNsuiL55ZTf+2c
uXU63OtT+DmRQARowcJHAwaZUZ6/voKiDL7zc2blGmxlDEPh8G2AbTZR8jYkjYlZY+lS6qZ7luYz
LYwIeehOaLBFWwjdD/xegyQ5XLm2EhKLRgVXiNlfBnPOWRpoJotnoKcTNy1dRycMcYpvpQ8climn
E4wrcWa1idVLRFDbKsfnQI0RgonafiwzBa3xU5faxX1JSWMjZYCe442tOT7p4/NYisYfvsZLcmGz
fyKJTH1GSjHzS9NmHikpjaQfvK+n0NjTQ8If/DC7HYxuqXrg6Y+PAwdQVxk8BcurIj46jOn+AU/8
odVBKtu+POWXDUZY5Xywbzc2hHRgKVIVhFP28EidwE9vS1MNV1Bj3R0aqKp8vSTg14bBT2hUZ5k+
DuM/axcmOhTE0AVyCQSXafUOCemDe+Xr32WJI4qx4IpUeWKybtSVoNgiYN4zZn3+06C9qoZslcGm
EXleWNh2iA1nGFdsC9ihVspANcppifkNl7VfOeYUlU/6+TWS5eIaPCuvpTMCRu9Awa5FvRzY5XtI
dDTJba1acelLyjOv9QNv/ELLNG5ioigTuPaJMddmtwnEPbB6qrLzRewID3/1YLUBd5s7xKm3lrZE
V/2PAe6aqLlfm6jJcsdAhX1mrOknddJlhzsi+AFgruuVpQbyEh+qZoD6a/QceWOwk0JYKspmpZ6e
aRZN8oINXBUiqiAUCtGe+yI0WOMD7LNQkMAztfPkVjCMVEGz4FDCW/qSW7n1vHG7foORwRIcTzQH
We0NTt3aUoGpurb1nC4b7PtByfuDI+k+hI2EKMhUC5sZ0FVPLQcTBInwLkkYbTadHghiPkQLNqxi
tnG6Je9ndQTa8j3t5T2nrl+pcLuJ4BuMIN0/0jiOK5szf4wjR/jwyukEBGZuK2kxH0e4OtCuE4Xe
LnSoQLNvD0Fb9RYVbyzz6VPNTUf5lkCgVPd9BzK9ENLFQ7EMaSepSJQDaM+amz1c+CjC9ypIem9j
FKeCsKu7nNqUXlL4N3KI42qJ+5+adQ3Oyk0dkb2bi5KXWl9UvNs9ju0pjiWW4ebUtRHNQQihzu+Z
f4gPkal655Wz21+bR4V5Yfg+WCiefC/mm7gG8SlxHD3ItsIcXwehOAcdNTSd5BbTsXuR1hMG0uRd
gkpXn4Bri8CnENRGbLrAChvG1Z6T3J/DYUjt/4hAnAgbJj/T0vwuEISyxug0HoIrFcpMuuv8OzGr
8phog81egG5WPtI/eGo32AWopO1qq7fp3E/8QoeSvq2lrlF+bdv0cAj286TZzAwzkK4dMRa0qo1s
uoyxJ65gEq9e021cL0926xGZyVUwSMM9UNrR9AqjVsSqGbJwJtU3b/5Z7w6VV6gDPS0hUdEOEE20
jxfDEgaDeMxzys6U2OHKVf7WxKe+3YWrqaKgU55MhbaHD1PMggt+EQAdJU7bQjdhcELOC7ldVSHN
+riVyQP7UshS/noeO3QlFz679BkCf88fL0O5lHVlSCGIBcGd/R5zcNeFQDdl8EAiFMIXbSXG7z/j
TKUXnmf7jtfEHREa+qrPYH1ziGQ3mspwsxH587Ft77+pE0POXRkWqwKdoO+jfRH29kwx4h4vW+Ev
lU6SoWmCVWt5/nDI4zmzcPyS89LbvEKAAf4RrAyO+GqHGPvQj4BkbfSA/MTFCdNDBvINeymvUXxn
/CDreaxn8qe2lmwBSjK0t0KjTw8EiASNrH5BiyNl1Q1c6PF5Nq486MXd8w9wYJmiWGC+BV/IwK+S
j8f46rwu5GZrvcVCgTQYr+zWBTgozNiMwKO24VpTBEZAbOwdTMScJfmRFi4uW2VzzBnzR0/fSxKQ
ByNgKXCwjxMgroagexozQ+TKo/Q2dvCwINWHOJsbQ0GH2PjegLLyz/GnXQ7hHlDYyOnQ5Tw+XE70
J4nX+7SrhpqsY5Al6gugGMhy6MyeAgeoNB4td3mtv0NyrrmElUmnUoesEPLQztofZs1TTGO+GShe
qzk+904MLmpt/2j3DlLX7nQV0h67AbZggdBRwli9MWcoUafnJWjBgIvjXuwqoUUxoN3AJhUbbT8d
9U7W+aK0lGtMitdC7iWIC6InSySS/HE/2vA7Hr8XFij/VikLaKhoKaHbadqoyfsuI15Tu8Q9GVjN
ozVkDem3e24eKDKNvEhBXLt7tPWrc96di3GSqI5gN3Z3o5L17HsjR+pWj70G2JBYW/p02+ZKjdDR
pffalUKG84ECIQRxfQmKetCrO6quTIjVy4HR2t3kjLUztPzqBC57vXGTDvVsLvHeDdHaQ9GLGD+q
0R1/rle7k1noZHOYxB51RaoYuIHRM2WmQGU1skHEQLGXy5stSDV+xgefhTPO4bdnNIaWmFltPzt1
J/Z3Gs6iG+mfUzB6PvMfwL5QJxil4UBNMZm0z1fl+D7xY4BA1MLmGJmOIF6y4terdy++hwyKjbBw
O7tA59ECvBwcfoqCbs3vucOmkYmf66a/EIwZOeLhbfNF69WR++gD5Funh3wyEixzpNK881W3T7sS
v8LscLF8cffibDHeBqsxITYWS8Sr3U/AaYWCNV24I7vQ7wb/bu+T5aNwpuupL/lI75UK3O3v7M9v
4xf3ERScWYIW6vZmXhTphSd0wtMdEQ9oNgUDkJSXSRo3nh0QKCH0KY7ob7iHCJef1sGrXvwMtZyA
4lsjdg/xASxsyazAkl48NJeW46ossOTD3wp4mui26w8DF/un8TQ6B5c2bCNV8fTW+FT7ukiP7UXl
CxDxkeB5X5PtFTTsxLGdn+ysH+aAXrrdlzGn1mRdqZ6UuazO5jGNak9H1ffzGXziQY5I8AsqGCRd
oKgrnp2EjtuGkX0xQrnL6EVIASA2nFKUJ78DF9zD49TfwsZiWrCuYgPNEtwrNeHhx79Q47iGaqal
e7vbkrX+gb5BGKDJr3W6iODDubGL2tenBVWnBQ7RTUVFBzIGDBbE3X6FwWM3EmIBoiREA/fFOxOJ
6prGFZ87r3U6ovnBJpQtdaLDZ/RB1UkAENqGaKt2vjiFbxnPQI7navIohszpsd2HwS4bf3S27EKE
Mcptr6oWf4RQpDyPVluM7Rbjmg3y8088FSyOMKngEAIQpRmd/xJiouLkqPt7v9dSM4WZhUocf4jR
U7nHbg6xy3qwlLLc8xUvRROjBswZRWhCpcA5MUQzAdn9KoXI7QK/ebDSc9tNtupYed3ReSq2mgMi
mKUhGRY87cI3jr7S+hHS2TAQTfnOMyKF/h4v95W/AO/os0UlnfHN6QcZ/96SXtb91qkTSKJvJ8L0
cwIJ8UMl8gNiEj88uOHX+BFlEJNBGw00B/QpztBEwiMhD+AzjNfyt1KwojO9KfwjUQyCQ/ZmFMd1
UKoxw5OUE1t7tTUrE3WE6nYYDKUxSLfJMhcVu9nen4vRQBl/WeehjgXdygkMge2iIgVWR/g0NVBM
jeZXeBaU+b1M0mlWQ3/AzepuIXsBeB0K8lec3NLW6o1GnxcPvyQ6/bhjxmPq3Ahu+U9Umey09oQT
smoeIrCFiAzUwTIg4/RnupugNwdONVTSBuvTDRnveYdNOUS4dKgyIbk+08Wamxk7gfEDYy9hGYHU
nUxl/hu/49I+Zhpu+sdrWHJIV0yi6SiNJOFirGJYupVLcawNGkoR2cD889PFBbGyR9MyF2+iAbkc
z8PWS2b5es3oFfMUE6TxZvT9ZGPuKijEMmwT+c8UD0vWlhfu91rjUdRWHoN4seiGJ5bGjFjHlBg3
dTjDQW07GqcFqYEmv06tV92G7lblK60cc6klEby5f5ua/eoSPlFUI4OzDEH8rV3s5coQdsqqfXiH
cEPDF1V35B7HX6+29wlKiphUkfP7M+aWmkOzj+YXpGuc3vNVqOCMK6vXGItxrfCbYVsDEVIPb2a8
Zklal9Z00PnBwnH2f35Hlth0V+zTIvde6QJAkE0kiuxDE7lHYYwkYblTza6RfK2VTCdCx5krxPLY
YMuFSYGa+TdO/ui/0i8ufU13mVtKtWUJYKmRiFKYiv86yS8lsHwGftecbrqjQ141qv4aeoonPK11
WzXTwmbuWPL99FiO/q9ESHP3KzNYS0yRCzUKGKn0uRfa9ag9Cg3XuIN7wfKd9m9sOACGnmPCryNE
ViDKhLsmWpgSPkdMvyIc9Sdz7iMYnLDQZBFKA5u7tzx4XAZ5TTVEEg9lPyzs5EZxKBya5rA1F6zm
iCPNXA8YpCMoTFv82MITDysy7oAM5Oceh8Ye/RztPaapY9biDw95P9PGPuFFVmmuonAPwe+VjTGI
/Zsr5DwbMBpZfAEBhe3ZIcIRmI0hjkw3pcDCRMkheodcFY3hKy4vCRgyZ5clQ6+r735KVU8rs46n
Zn6xO/PyVWP/WPItr39c9/fp+R4wJpuOpj+vO1PlfKWEx9KW3e0VRPX4aQ1inkqKf+jl3MdP6RPq
hgGBimpMtOQ5cgsKkABePQeUekXo7a4fDSjzF01SM5Wx7z3Nz3yAin3etK/o3nH5J5rztB2iXVVN
a8y67+ZfqjlyOMIuBJGbrh6+vrhMx/m8aRyhBy0oUEvO9+hX8FHPqPWbU6hP9aBwPGBAFZB4oLxK
yv7sqKtrstTh0oiPgXyeENuVy3BHRDUYl1k1tc+fki2/FwNdV2Em08lcXNPyMiwhgRhxR1mmhp3/
9KoRmoO+tfeKBa8RuZaTRLi7PJkjE4w6gZ//cHEByaQjQpXNERW8Htalrjqk9Fy28KWQhAn0/C8Y
A/EX5wYzl4EftV3ztx2OHX1rbzgC6svGtrwdKqQgjfFaRVZSJ9om1svzjaVeejSqTvjzDaQU3Lc1
GP/mldjsVcH7nhWoe9oId3SMlQicvpcdCvunB8tdW3/7jjS9ywbze0YdE6c0R/uUZL/ArfkwoYS2
Mu0e7nvws6mQS42ep00A5fWxM9xMk3NOh2NQri0bAceP3QvQmhC1wfynDkBst1txVet+eytUOX88
JpuVN7/fnokXnoVax07KML+P5HRJ8cgPlVHZx27d4l9w/QoF6p89yNBQVV4FZzgyx0hv1AyqNhhy
TT0ovkNetQDuDvsW8Kt1lmyuWno72b6X8ltPuxbqbxHgt7gkS0WFa/DfHwNs0h4fy6J8WOswKfRr
TS20BV94VFUz+bZXobcbwdr1dAdEUZuQDZmNlUOpffEsCNxOFkoW6Cj4EY00xlQbNVtaKOaKPcsq
bIG71nw2mg6XZ4TglSWi6MRqCrbZkgvHBjzfBgSoafcIEmyujOkI1kfvaSq4RYEnzon7Duyca/lS
Rapl4xkb4SdGeDMcDjk8TdwlB1jlqCX5S9diukhm/D2rbkcj/sDijg/v8G3dtLRVBkzg7KqD2iUa
8p0nxqf/XbhE1HYgJ6+fUBDy2L1DNH0O6qJ4rvIgaaDFXweMTqdJSJS9KlFmTo8ZuSYDd0OeEUbk
REqFVud2RyCzVjnGPC1bqDTiN1RIzB7LH4/1zjB9+mTeoV7jkOnZIFk229qqWwmxW6q42mgRJo0g
uqhFKuCj8U40woNMwUqZGxP7MQWd47Fy2Cu7slzfwaOkV8QFjDksinDoctZ36D3HAwNQNq8IQkHR
BAAxltzDaQmhYGvJUm4V2fBv7CZLsfPOgxTLE5/nLKqyQw2KnoY/6r4X4W5zG6i04bEfWS3EYS5c
unUOQRHRt4xzYYmSvoTB/9uY/55WR+D69JjFbsoJy0AmhnAYihz1Qjwsz7QkYNNUDmT7l/Qdg8Vd
NBSdJWErwtLlLgMTJxhlDgI3JlhO+T/LJ0vQQ+i4lqCF68uxtgtPK65qH7+Y9soy7/VzL35lz5jc
T25Sj1ymcFk3RC3MT2zT9Aj6Q7vSKUqRRU72gYQ5SndToT5bMRSAcMk/mn5GvyLcSZRoOEEX5zok
mmS9hT9BRYQ2E7pTGqxwfzOhSvWYv3s359FQfVAwxsi6wCjLzuwyAvykLEn8MNtpzZ4azPdz0nFy
W2zki5VEv7ETIkW93c0Np0OLqXp9zJi3CF441p7NkaERnUmjqNTPG3l9l4nCP8BlMtiYyDAlUm3S
wk/WSCiyrCqtzsvLMUxN2oMHUugo6xPm/uADqKwEO++RBTZadC6XQ+OWRuKF4vkvV8iUW5EN0RKk
lXQDQ2MiT+gBvwMYqIMo8pU92hh1Dc5oxP9T7NIEj5IhKIHaNmedXRiBzU9//8F2QD/katClA/FU
tQux+r/YWntnk1RngXLAatWzjLsYTJAL9ZbSSecCyOq9vZnVsxBym1RNMldZgwrgkpikIIl+2sBM
y1pDTVF0IcoB+N2WEoisnePw1c6P8/KWZ/z7RFwKwIBzzMfVtDqaBXRAS5j6XiRxh35YtLXoPDZx
jgVEZxw7t4qO+eUVM4mB3y/1y2A4BXWe5KgbmXNU0hGEglOzYEaip6PBOOLPdYdbTAPrJNwzQoKd
qbg7d/TcJhzxxdx5vvcvLms7hRxF1he1CESXnvSuPgbnwYFckSYcFg/Tslsg4oV8MXF6ciKx6PoT
IZdX4EWWnhdSxysFWUteCofIOiyMDHmIlEfjOZoXAaCeFMb+7U9FWz7dgbNcm5/21EaIk3xrjFou
cNlCmqmIee8LcivEG362/Emth3v2h2L+Qj1IsV1/0Qve9NjCiPn6pqzUUyGUah6BwqObYPakbAQP
CchdEA54DvcfSklBpiFbs3701FpBwa2o3ERhToDeTwhDzRKT7mj3gTHFoG0YPbkUGq6gzBgot+1x
yQoxnq8HG9vH4DDqg1QbNrJgelk1Obfn21Nm3k8mT3zAiHteokG8SPUz+k/u4QT/p/L8ENRiwhT8
fkQrHQl8704jciCN7AylzhQCNofXquLKShnJo1da9wQOfwOvcsJljblay25QhR3Z+ZbmKmu5Yw7/
g7dbYCR5DBD3H/BxStDhc8eTXrzpvofGmCXowevRTjJq+u7s9voRb1JoSWHoxMj4pnjavLBHKXZr
SnqXX/+MFc/SV/On/dv1zyccKc66nbhFApD4QXzRk1TDJyHVot15eO+kOy+q/Z60Pzw8esSFdfvf
MphghknfyynDwNCDVwcdCaiWMueBQFeuHjndnmtevcO+4jm6fs7y6k65vv8kFBHy4PfpzDlk9nlI
5O+SdGl+TI9wdhOSW3VKsJIDyGPvOZpUcWHi0hIzs3M3qhRxLLE4TI6mqGwKUgM/hUfixd2R9Ly4
BCk2Li+hoi4tATloCnLgzWcOhmXPf6qdQ8t6fGBFwQZj9as4wKuqjw48Y3M75EXF8q+olVcPmqRo
6TqCtdrSv3SNif/Er/dp/a8a69EXJfF/YrnbegJg4Wja0p6v/jcnexoxh3w6ySqbODDCFkvNfdFG
EjPhrMnNAPOITR/Gs6ryaMip7yN8Suum1V8CZ7z1+xM6pzpDsQVjcPa0d9HsdJqHksQtxQQfAKcx
go+JYiszLQsqn7R/lDKyuxRVKfwIpd/Jovs/ZjnfZ22Uy31GhQfShZ2iA5TQ9vhGHZoSqJ7NvZI9
7RSl9vJkl/PIhQJtJulUxKM1/Si7KcoKQml/An49C/4P+HTVbZLhQo2YXQftFzV5n5394evzvAD4
99X2wBdg29POw/e+Vn+VUkfjOKedrXQkDXv4SXfPgb2fq4oATeKsq0mN4o21pmCO1zdEOZdNsiKA
AtNoGpEAQwzwRnFJx15+s3WSVMKDP1w6/fj0GiHKmks/Q4EY+xVKaCJOI3tOWObErpIuBaei3Bo+
knMMOJOTO+9hMgG02B9y8HxsP1f9686dyg7RE/692L3Hs+fFqvL84t0dqFGV1sxDaSOtsAlZuNNa
AbT3wLMlJO+70CuWSDEdbFjOCCfwxKQRt7usQKB55ax7T2SXO8tzvf9XDBJRn8kL4Hkdreqzq5xS
NIRhnzEYYz65Udo6OJjJVP5xLLZAZipoA0gXIBcVQnZN9X0SZaaMxtgpeLP8xnRTBhIyPDKGSESW
NZkolzRdmDNdpfpgaYBfH61SPmkhqogUc6SuyoQVW7tSlsBEg8YEsbVE+6SgoiHLx1scHFBVfW6R
5vXV+xfmuiZgM1FBYFmaI5cdd6chQLUSJI7pzvackyF4vA++R5+NhKmDaOPJ65YF3FrChWlLTo11
BtpXJ9HdB0ZKwst0W2rFJNlH9G1qdoBtTb7pF82ry9QbuEI8DQulKGn3N8TLPDqnFx6WfUdmHi1V
RtCUGO3qSioP5Ih2iKens2ukRSvHxd+JOVmf5IYF12mB9lVCGJdpgAaOidb2FpAdBsfQHMzA0IDi
ZJjTe+nVRuVjgUTQDnw4UcF7XWPDTD5cc4WDENaKFCfU/Bf3T2wFcRBQjwjtdvUZ/PC68yKcbCOT
t4CvSeZmby/r6KjeUTBNJ1PuwB2Cpq3vlBskBvfgjeLO7SZCMXcRjRniNBYDUGbYgbQSfuNxM4ZK
TpAgzdEGP3xWPrkbwohBPgQfOfoHxTCm9GgVR8zpNi6cBJQgDRpL/hhyvzM8o5I7g7J5LkM+pylQ
Pi0UbftWHeI3BUjMhnVqIH5N9Ibc9hO47AyX+Vqn24ysKmAeRCL+YW6iBlYArGK1yF3Ik0JNcfBy
farP5FwfLZcBDc+6tT6XIVfBZ0Tygb05oaN4EjKCHut51M6+KB9nuvQsYjdjaaZ/FZa/WlsJ8JXF
p8yDTadmhbdfFWCQ1tPhe08b2SEfdZfOsl++iSiV7M6Zmj5W7oyOyqbt/ss+pE84ERhLdiCby6ec
jYGoYohaLigLw2itwvD9pIag8J7BbILuHI0uRhQ5Ud4EUKENuJMdVQwhr6X1lae90eUeoG2HoVgq
jFifXbd0MZCkzBAA+TWDPws38Vakx7aA+q2bY+A4bUrTMQja404m2vj/2x2DsQ4eIPt7GIbg9/cY
qYIJSl42qF9qaE1DON4a/Mfhd4nssVQyeVXlIMNqk46ZC/pm3785OtKUhzu/z/3FIClUpj+frIWg
uJRXiiTKgpgWItFHLYoBDsWtmMZ2gCVUZ8XZcTxguiS2dpZ4025BGOmXcAgcu1Tfb9jQi1CcV4n8
Li/ztf5yey+Yjkwes0TUyt6bA1vxl6Df0Lx93j/8Orr3UZ3kwhNnW7lomHReuhPEZnFawGxDc2do
Us53e6Tt+fmTSmg5sJLxLcvgE4g0jYawp7YaGji0FpAaH+MiyZCKDztN0WMy1KNH1m/AZQCNmc4K
fK7n7pcNXXZxsNd5DwmT90Ij0qGVbztM8mzPZiLJM2oZkXfxWmqx2EkR25/k6sRVsuaKQ1TbNpYy
2yxFjPAmhFAf2zHwXYy0nNq3qklcJHZp3Tt56GKGD1hbdLnTskvjYGs0vF5QX2+/LGhyhKAjOK90
DK4LDJbe6xlzhHkbZog/Vps72rRlFXrU2//WOEtRPnGscj31qN0+kHuN5Mx+GtptoxtnpnGPbHC0
ZOSB+r/X0W+XJO3q7l3IsNfPC1OiTHQt4y4IpQpLxX+lvNw0xcKHaEd8rFsPRkY9m6gXyUN4MCM0
mt4R3TbwbVIi8YNrOhBtDbQZyGsynBnocuinHr+/IuNDwkVAeFzO5t5FB3ahozC+mFzoqeDwaXzg
18xcCoW7TDfS+Qq3mv4kiuP/KJVEs7TbzV3d9as4bjomtH8OkOEh+LpQVl2271/Z1d0QPO3xmu6y
/JMECpoytHnLrVe3dUS6MN0xbMfxPbijKRZH2Ve/YI5X2s8R0n6a/j66KfolyKdXDVAi2TCXEsOB
Hulf3y478GHdn2IrE7/N6P/VUpF1HNV1ZAFQnSbw0DWzt4UCwSl/UW/1MOcMdy5HL5PBIPSLDDXu
ESymwZ0RbFXMUkFLwuS269ct/jkYANF5WqSwKPcBhAhrewz64TfpoiWeGJNg8W//apKlc8Cmc1hl
PSpllZxhdKFuxxjL0RQwPZ0FyShUzpWSQnY3Q1IKT/5l2jOfEFHekRdojf/Gdymjaa6+/JUNJDd4
SZiUeUIWA9oHk2Dj4Ey3THTd80DwfYaqTpZJasS5tlqC9vcsP7OrQs8bEMyqcCqTzqOrCgTEyjoA
XIoaS+2ihMFbRHTr9WGQnCUn7qwHGSfXwHZL+LbwQvyTOtKRN82IzrGNicbGru9aM3Ntu79jAoDL
0sgS5cLN9sH9qdNXMj92d0qvp93RXoQvVTkzOXxcLog=
`pragma protect end_protected

