`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ZP5ShdLS0KtzNPc3+HnteH8XiWJnjr4o/rZjRqBo09OIqK2WMiWOqoqyCwhZzg1fmUBw3nvOtnGe
5KN31K6vhRFDueoXOLv3kjfzeyMvvthDVw20E6YNN2El73l1nIM7gI0zZyCbahxou1QQipebJYSo
ohh6Ar1WUQVr3MUF5ZabbEtZJ9OzMibkfwx7XxD7tccOrUniMviCcfRLM3MwpBGhoEjYvB6QnvJR
KtBuXIkDtoXndQXWHyyzrduJPOKjj4FDswaSkwoRQutjvVaDNj5t0xYTVmJbD2q4/CzUibWy8Tdf
goasiFfFQuGf4zvg5JwL5DMlZ2i4GcDfsMQ42w==
`pragma protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
hV3DUtdjh5cCXhAydIygfW7Aea1WD7msmhG/ESfj33P+KxvMQO6/F22+fNqhRbFt2M8LZNOKLJIW
G7mu4k3rmbRe5yPZ2mPShrhwYg+HS3ZqaoTGxM1LJk1aYm9NBpcRs1WHasI/8MH3h7CcMm0gJI1n
mhtMKclIs5/6jC1M4sp3rt4y80czAvqoWeA/z3UHBNOWSF5kJQEjunMSHyjz+vV4Ex1DMLrLYI7H
OJ4aLr3c70bC6WunI4cOXunxZxVqxbU8OD+UkxrGX2+SpmDcN8+EHVG2o+kpWZw6dsVyVnZ+SDbw
KyFl5jXQxPDrI6du/D7v5p/nsW2d9ma03qwhXA==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
PCkCV/RHcI4lAdwSzbQFsa0gc/Fl5SDTI02JKr8mM77cJLOXdTRM5Lpy/NSYNrXCS78HrDU/u0BD
+JHuBrNvZA==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
fsDa0nx7tIAwD1ymg7EXLAbv3PFx7wkgwUyft9XmJ3K+E/bARUBBXp5b6sUDJdO28EJ+DPepqOUk
NJU1EEMf3il1uP1jaxZMURRSF8xRfhhMyt9Nw1bW61pVuRAZyHcjmrJOqYH9LcLsPWSt4QanX6us
KYLjV3NTodhnKI8A34jtC4o+MZE2yUrVPI57+4Edl4sPOuJ+D6M8S/MA5pHQksftxAD0kAbSIexB
D/IphNxyxrlvHHZvakCjMZFBivGJPJrBplF7oMrf0srfMD3W/+6Ad3mukPPL8Zu7zT3bRO1E9qxe
+jWLo0L3l7AJOePt53ZL9Q8IYXgc3W2uDQE37A==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
SwBqa8D9MuZaAdD25Ohyj4f75J0CK19aZRVLA6+npEhNilMSaDqzKiQEY8KzcZ47Be8y2OeAJlKm
JUBjYzuq1b2fKY/DmfeyPUmHs6LBmez9s/3OlfimLs/08PJC1mXK4zcxjbOPX/1r0UReV57qOlV4
k76a4U1EBC276bgklYk=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nncslmlGKpDTG96HJl6inWWrb8hHUB3OTqM9lGYKFy7L0t+6a49M/T8FLOL7FHMTpjS6wzYdZWkt
EwHX6jOEnebNx7eBUsk/U3PXJq/4hswHqvDIawjMpwmLZMH6kSgrnoO3yqAMRJNrR89/oQM1RyaO
cbniWHQuVLYRLqFHJ+2na2mz5QHpIyZIhMicFrEpNGuAHRzJUUc+Oig8eSW/aTsuWBdntVhOOEFW
3fA1+yQmUWXoawoIbo2cjqhH8ES2wd/BWP+YbW4nGOP1o20fOU4+C4/Yj5dzD7konYZuhwfD4dS2
Vpb//CcShSawP4z/9VIz3xxd53Uzeuk6pLYO7Q==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
fGsyZLTlW4WCvuwoh7rO+ZYK8cgUbUlnS1MyKsFZZnGX2W21NiXQxymtOe6KM7Q1NUe7r1vR1J6X
CBNNf3NHI8UPt2KcBs+z7wc3ITQIdOUYw6yTtUUVakWZ2Q4Va8mlKXLD6w/6DkToKovRvqOnu/Kw
flQOuJ7DTIuGY6iMzVparpNHVOzK/YswFZCHVcdxdiZ7vcovzKXMtVRj0y858wcIJ1JuXwq+oT4a
lXYXO2MxYfmgI56KVd7g9yjg+Wj/RUXTsXPmCCKTmD/b2STBmOxx0OTwBayli1lLNS6A4eqIv/bv
EHVGK7WamOBTB3GYjJK2TGkocUxdIgklX7kP5w==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
SryJIdaHsTXUbI+ZZG7ntJU0Bea9qvBVtG3mAgYTGHUGj3AVC1WfDqSBU2dD4bBDWBLv0PFAfvdR
oMifCXkuqE4xiHpar8FC+TLZqM6yFLTPS3eCPmp6orz+Z5pscy7zSZLN4YE63CxNqlHRRNHvaA96
mQE3ULGUEVQP7IVdLjg=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
DYBB8c6dExJlWVlDUSBnllEo/IvUYp+IvkcLh1lr2QWVv23NXgdgKS4Px0x4CpFpTLXRsGRY2/iC
YEvSLIEbU4DlBKFPZzmW5aLlR6BacF17T+vnxsRansn01dW+aZYn2QngM9YxnomRUpVIuzkaYLtF
kWoRSM/DyXvOzivoWKLb84FkRaJXnnd7Wl3H94o+qLR9g90KU9qcRNYBaJnwteik6AMZa3qF68bN
VbW1pdUYmGBG8Yn7omNqIPKKXnmnGl1R8vtLPdptz/Ht6nae/uQtkIMvMoqW3TdO/79GO7tdRixb
F8dWR6taXuLsckyt0txR4M2ZPqdEhjskOezssw==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15424)
`pragma protect data_block
3uZ1llwxzhDoaFyACujmlhAC1ay00pU/050AsRHVZh/9atO/BJ+03N6dnL8AkTnDDL1hMfrDNzYs
tWp4pQEMh9NfqadK4r6sqWgBKta3MkzRiJSufoLmRNgbV4g7j/szRQcAeCz1Hqi2GJtshqV3gQf/
W1sy9xqQpUyy+K1ouR2ynAnKxpX7Gkwx3jSAV3HNYRZUHF4PGHwR4OCi52B1az/43kHW2cqR3liH
oP8xUKV2PU+oKDfhKL/9lh2RZuOOzgBs86FzCnLZ7AFoU99MFXyplH8C602yh5dAdfqUAheU6Xlx
mtH8UuUUyx/oJIlQHYvb0gozyrO83orAgX5IV9KZxZGABIs6ZQgwB57KQ8VPhHrIMTvWh5QTp0PU
dgPM1sdfkwGL2r4KX6DpfZb4Re0/A6v5Df+55WrF69jUPAnIIB5RuRGU+kEnabTQqAz5OHLMcOyD
cYPRCpHrDOUeJ54LqPACUMBJfGMKy3cQx9YuTxAYKTqN+ObzxnNa9NgnCwMmkclUlOtIBhIALSvH
eXPMpC6FMxlt9f5VgMkxqI5y14s45Lfh4D+nX5DJHU4c4E0mbnOohqyUJVA6zUzxyQotbO/AkC5g
kr77ES/dqoI4VgWAoH4AYPlFlBm5ZfSm51kbacSh/0MXLKcUE6ZczwbFH650LVs993Dm7BjEhjcN
7xUzXy75yFP0BXTzlbgmpyEyYQLvvtNGTMw/WVXPAkCARmI5n5U7oy2eJLQFoTmvoSodxsUF4fQ6
+MOlyBjqF7s1iBoFfyWmLyMf0cSiTvLtbOg5N6p1b+x9CbUELuleXUWAiFhxYGkR2ozyCFBOezeU
2rmRR4uiJC0Nms1ZTdvdANdh3QgGFLQSm//9OKexy3FpOVev89IKQCLNYsM71N9A0gR1MibjONSH
Q1no4NUsnLYM6IjaJmJjGR/e2KIklyAth+KGpp2S4QK+/Pzi0xmZMNbLEPs+DCRmLzupkC5JZAYZ
DgktaFTLXHEKkRPsG/iY309A8Ch8FNrLws9XNHQHDWZSGa1PSk9zRDNw35oPX/WR7PggfLWwcIfd
beL/oCPLEJ9i9rcAL5RkXVG6DL+lXhaTiKSLxngMXVGfiu2RpB6Xwe3QF8ncBpyHb81mZcl2lNvA
H1YmGYkW3OKKBoBJX37s0EBUZvW2WzG+Ugh/sW947LIOuQAlSgvay51BbQxnN00y/l7RpfD7BbSy
g87iLm2DU5rrfd5ubo5Eqwgfqthsj67K4SY8eqvPDyaL3hQe7g8ce9ok2g11p53Ge1uBQGehRzZ9
s9HWoaXcGZnPHgJrCWtD9MNRZapdlVUSZUgcKN8m1KrDf8tPjJaoStOGmKuJ9VZ5KuZ9+u7gy6PP
TKPmpjedK9/g/xWyCYUB6NxxgdtS/BBi9G6PDcZVwR0wKQQdJZG2/1DBpOvxgS2uRyDiJ95PgQ0O
Sl1QrVDXc9iUGmrg0IYtdOntJtDIreydMek0YxuCKf+bC1zi/zuTdd4EVV3zNhP4x6DoYLLiA/lA
wiVMMjSLlTl0j2SXNcAMuWlOx3zb0/3oY4trU6pZdvm0fNnII5ctUPMCP1tYBWbxItuhP0yIyzcQ
Di34ifjJ58C8F4qEz1d9v1JQhi5OWDbxZgmMLw7oxIYUAfiXgnUFHcOY2GKLSYVjylNGjXM9Ihx9
ja3bWPB7Wpc9wra4p+pdpdy0kRP75zUwjUKUt9wqPPPzdu/VnPhQRSWcfZoePsSTuVIp1coiRkn9
NHLCKa/m16Th3cAP86GdqF/OI9KJEtCquQkWDs1x7PEuKujb4QkXASRjWS7fkO7vSvWSVJv5X/r7
t6R29Cdz81KnZkVTQE2Y/eLy15VYJ5k4Uyuy/R+GDBWWoa+6UNbU2GnQXnOVn/rV8yzhk8M8LfDD
EDhMKV7wiHddWwphtd7Pf3wHD7aZh22mQmDstPv5RvaeePYm8FoKU/kjl+kURcHTrjuDkvEo0Pni
bF8cNPad1wquYxrENk+NrWRfDUaH+saQIqVCEFdJazwppw47n8Nn4bZQxYujRkchpDFV4FJJG5jp
ac9/khgboGB7C6vG5naBRBqDiDvIjwVkdZaZMpjEqO70RChCV5NjPuNZWozbWI5zJ9ms5a+Zzngn
/OVYi0saHR/FH5IN4wzWlSB8A0eH6S9wQdPoUnADb0ZheJTw+HoO2e4l6wcn6d/XoDZTbqGc6O7P
kqNklfSnblQdKasW0i+qCy1DqSW3at27vAabitHPHYFTMu4NqxG3siXu5tY/M0wVhNiKMHg2lY55
TzaueFQwnYujToG8m33TCzsAf4ybVuihyXXFiEgvV1KPjxXG2DWoqIRJA26jfULvYoZDD8WUxKOw
LtFssZ9x8Do+mU1QYLK1zd9WIfuAvswbwy9GDYJsC83iurnZuCXtMgwHYOXquru3dP4FLs9NjY2H
ZdO1gzfHxA6qi02jtUgX5qcZt3Ns3+r/MQVRwf22qrZR4zCSM4WhWB4Wp5gdJw/SlfkO78FpkmIX
Q1Lgkh4ehbvl2WHBSSim6NHCTATm5swy4An+PN117D0izmqEwyVkzrjJgJYelqazNo9Ghq6g30U3
d/sRtltvLFE6NIdMPPrhXvf+fne3Pw59ofBN1dRqJEZs+FfdnHaU/NxV0jaxDJO0+pzWQ58cZYy7
W10CIQMjhDbHqqiGjJervSH/LNcys0n0aH0bqj93nu5AjwsgoH2/b7Scc4MQHe/319NPA1zRoZpT
GGPTvRGKd1ZhWfj+qdXk1ctszmwMWotceSjXvf7hafkbq8VSzHPPwUtdCbFYdSTgH4OjvQNROvWF
sC7Qz+6Cbib5qtMtNLDQtN/6Fg1O+CmJ20cszqv+HmUZUP2L1wb/cA7KqQ+D3ev130C30ZzQeTr/
GigvDShKCpv3LN3lJc5V1QHhTQMhP/AsSSGsXl4ls6Y7GOZkjGiv5GxcAX4NiJxyHJ3++WtmuVnn
HWPF07zYKD5gsOKRIYH+NWduNJYp1kAK/6V+O4XAe92LMu2yqcOKh8LNFQ/vA46+NTFUGZkUJN/x
gfCfj7ilh0lRl+1XdwBlxpJN4KOtXXFplmKzZ5F2RNrEu521NTtrQvqbWfhEiE536QgwYM17J2gN
oNZqVkjjW8AFjsUzmBgJKo9jh+iTSbyAR5tbgn6G2xwhqZGTxHOSZpg93H/Quj/FVSaIrsRhCg+j
Btao9pEsm+K2E0OWEq7TPFXyb2TMGLnh9c2vQytS3p7ip2YHw98uH4eCo5MuXPKdWut29mz8Rta+
5z5afpp24fm5XhjioCGVeZ0/uirJMSN6J6ICoC7w8X7HTKmtkaX386IohtO/t5HIm7MKCR+eOWCD
0OtJ0v8sk+UJIGLdE31e4Q5a61k6AunUacVPe8kLNkzJqcne+R80oAi2NvtiekWI4DXNYxnUTvxs
BuY4O0Il/ta/cw4NsgY3x8qPUDs0nLCbMwRaibdAsOIIyOl5K5IhUt2ixezKKRi6SPi0H4CRZy4E
0C1ndD4phEzRRZJZPGQJsAqSv7U3M+YOBNGBBcfeji67aZaIrMN9v1DsgMGp6wD9QHO87VSsZ4bu
xDEhS4bqhGk0aCyIiNADvh4W2I4TTjoJED9BxMWkYmrbJjgRYqaaiL+Wh2A+3XHSd4Ib7aQZi7Ki
Jq/xgteqcql4Un5v0Xf6m9YXswOlxsYHwCUEmt+kfxx7TSm2kY+wrq93SPsMTyKP6WiUue0pXZES
6AZa3cCEk0Zs0FAa9yBTTKdR9zl3MA4krJMSIGOiusCDAbetHEGrMeNkDzTZuw0+vBt+gm+pg2oj
TiLclqMQJgCrFH+eOrCRd6t8YWfkUcy1S3dvvwcjZfSGtLn2WChSHSxWT184TgstV1085lzR5WMK
jOeViVuRd+j70/2eZpYuZsmGCvkyCgB9u0hh9PR5hDBoLjaEg+27JlQp6YJmzPAjYlp0zR7TBqpY
cEVuvfgHQyIKVyhE+QkgfJpRd42p8kWwgIjb8Sr1IMWbP5rCKgAZiLVWtT1a4cYSazkaOn5ZNFhi
u06260zXb6kB6zafye+NeAltA7h8mN1Q0Met6K5sGqyG75pyrk7QKwgBbtPNzNUNcm9rLAaxHVvc
O1T0gdvg7n5HOB75rgWJHLWZ37euS30TxcC3nONmmhsQcJWHhH1wszNEktU9sRBRTnJ3bS2K0SYj
jXAalzjt5PRAyB0/fPzzSc8UPkTAItQbEDJnLfOtYQxGo8/6NrO0ezQn0EDiFh5jG9tawJbL6OtW
mal+5FI9GceRaoJbCv0M5m9gfzYlO38UGIoY5Quj5uStMzty9TSyTLz0DSNY/Vv+F+g0ap52DABc
lAY/AFrCSPGPfaL+xds1fOT2dmX7dU0iLM90weaidP7OyDafUhFMb1BRDy0A143bvi30DbTJl3pP
PoAUj90V7J2n3oKat5YVzyABo050BYlbvayTnHZrmLFHcrbw9AC0Jfbh4fs/6i+dITnEfV7nJXNY
koShdf0PDlNzHI7uZps8bmTISjPRDsldY5FGBAPvvJUICbTNEB3LWG+LgxUpz80qLsaWojbcr/Ql
F7VIXPooSTtZLGHKHF6P0gwbge/wp9D11VhU50ncdfPKaDI8U9+b7EwDHyGjMqQZ42cwKFv2tBJe
LC7WY1eiygBGlzRyGyLrzH7qCuvxY2rzFIBrDYNqDaBXptv82tyHMI99egzlAr0SFOkXBZdNEVKA
/MQk6sGnfwXQBgzILpt/ZP6MdduGRIDCLxKLXBMSK3WfFR1oB6trlTLv9/qdOeHpdb/idtphTe+0
LH2/aXWZnUQJAuc6lRgMp8a9pKL4t0Kxcyip6vxzMUV7hzTYpqEbr/OlkuHSPideJzcKj/Ko1baB
IjNIKyoHTkc6nRS5sJum3KMfBhoxSFr2rslmcol8M9qBwALDBfwBwpdVB7kUCFPxhdZv3XDwYUak
lz6XVGn2LwNfldcqYN/HJmgDXkOGpW8w8vhtUlQyciuRpXrTzJ//dadhB4nFmLi13IxWnDIpmFf2
BmtVAD/ZdI4ck2JTreTz8Lr9kR8ymripeUcshHarxsLCAybfE8UpL2/RqiKDT7fKzTEmM/lShNQJ
GKpl41KkuW5OdKHXkdNZofBwN0tirVydgFHFqc1D9Pt7w1/BwO3aoqSnIJ5zd3/CDYmZKWPWapcX
F0TuC7YrvGtYIrkL6ah89xPmVFGMEgPh13t9LFR7pgKPCWluKem91akzM2iOqzv7jD47HLvY8yLB
VvvP8zIVLqraVRFmpLD9tjKqezFw2dtVo2l2G7OxpnDiI35vYLvkgTh1NZkMvSVyJavlYt+UfERr
7wAgncoWaOXqIxf+/PBoIEuQ1Ep3YOIJtXQvkSXV12YSDneCmYFYYwXz4/tTJoTjSj0840WcwwjG
F3Tj+fDREDTWeY2zUlugCl7SU3BXTlvysC6XqpV6hGvylGQRXIujt5HhHNhasdG37moUrjehif+V
KUgB2Y0rQvxz1WHnCaGSVrNlhNUarUX5AP83WPW+TWNOGSMZQdNeC2PJAHSKLFVXOljbF0XAxZOs
2GEwZgD8J6h+/gWrBhj6DuaM0FyBsEdFXcflPtuHdNEL6a2cR3u0G3J4ZkCHaVMAgiD+5U+yr7fo
h/Aawv4zJNvwegHt0tXfcomFyt2ERx2FJoZcu4KGyRM2LrFmr/7kv07HNrLz30FgaJ+Ty+dRSSni
YS5P11ttt466CbltGkj8NSKkG4C6T6CdGNeOmYgX4ehWdcwg+kQtlxtqvbj+p+6hQBBytTKXO1yo
dB5n0WDrzwlboEmfu9Vh3FlXe9en3pYZSqaxRl2+cpzXYYXacS3YGhHDoVvsS7YUHWj8hN+941Zb
p9YNdzORJedSh6b9axSjWRau1mHK0TYCuyIlnU766XbeRKRHCITKy1S3t9RxaL2NdTxsuDOZykbB
PVU5HwjIV53qfOQgRKvK+BUEO4Q7BXWnbf3uXI9h/woQoI9FOG1jfnpXw9H9rYCiu7oI+3UPnbJf
iRdj/06jeo5k6xghXo5sx7ZsNeNFczPbACp9R8ONoo+eEfBCy79gzBY68kYqyj20AZeBBhCepIZx
61MEKeMhXDOf++CW6nIKeFmIgtUKlpeuvUaVa7/R7ebfrkBRcJ1u6t3Lxg/JQgIcJ+JE6rSh+N74
rzRX0PCBsgIixaCtnHxLqsu46wLBFfxKSBfDf9yqLVnJ37N2jDcN9YsUY5UGiQFaSvXb1R8p7BD0
Lew1owGuXfR/VqXT+snBuDdFesUCH4tEKZXD/UAiI+XSSjxUVm5PKS8kpKDUhG/Aap7b/vc8Z639
S9Kfjj4WTsFCvxnf7BxFRAHaiisGLXn7OgRc4tzx+vzOaqHSSTzJjPt5wJjOKPVAQ5OnLyeppuvJ
RZPR9Ghs/lScm1tPksRv02wAWRDvUubrWgNFbRFjobhywNK1zR4vF0m3Nh7dimumtE7bWqtAXU9a
fWq9zt/Cy8Sdojqw/YqVTITVegZlvFtghqrtilb54AsImDWNklntd8Y6Vw3wMprBY+g2Dz0l6tDk
Z7ZXGpE/+cjlxzzTF9rXlXx5nHenMQn207zZ+URbD41QXxWs+/Vf1V/XfT42bsv4rdV6pquZ39Ek
1Zd3lZ93QdzN18p05ctNlSQwAZ9CjhA3ZuTwqDa1yEpJlBHsjEX0CBwiW0yWJNjYV6oVVbh3rq/d
BLvAlG4/6HS+TC9NVZs/BH4XiWy0WbYXqnR8pObCbiI2modR9DvlenFkwnSwmc61rf6wVUqJXJ9o
kCoMyK7C9tVSJus3yVMj887iTF0IrZzA6DxW2h8zXxV5nyUtSf+znFuHRvMl0vtA2Fyo4DB+MD7g
dyYJIqSivko3cvdPVOqeB3tF4nVACJqfapUkmQOsH09MRtGLp3+8hm8aMRalVRspicJyCDKU5GeF
PHEboZ1seXDQhKh08ELrngfdS+omHQ0kiDYUZau/gcIf8MGgaVgMyiAn4ISAA359wVW+DvBvsKxt
Lt7NBHHQrxQDX19mtNdraoy/bH3diFb/iPkTuqwbnbAgi721uT2Q/G/GBDCnYMGQwSNuSzO8CKpu
I+m1TGU6Jtl6xCVgJeR6k2zBBPsRlts+lbGreKZuK4/DJUvzdmDVE4CLPSu26wolPuYswLdXXPhJ
T+DZOoN3OcvVUMMOOEwysU8jasEwTUSHc0Otg4YAuMl8XEHZ3HvB75lEsO4bkB1ejfXCk7xGoWkG
bJ7a2ZIJlyenpwhKPcZvBB30MfVBfP61kdx/LwG799q1K1naq4FXdf7/jIXO8EXfBMVgALDkU0uh
0dciEYc43s/zn2GY3eTCHVaDWOZaNr7w8bSpasXDGuGGZvBKeLrsH1xDdh7cqaa9hoZtqbI75fqI
y8Q7KPwIxLrX60DfHbShnuRqsf2OwvOtfth2jF+GQtf/7cN284U9WeUeUcFO/MDod1zLd22b2fup
LBKFxx+7MHzLfe4KuxlDxU2ppMHSTXOVSyJRh0XreuEWBgh3Dd/p6Koiao8mSU2R+w5sDB9DkZz+
8J5zq12b+zR9aBrRdWM7WUcU5QALHW43Fqu+NcHafV2f8fO05encJrOqSl6BfvD7DSzOJl6SPHc7
Ai0c4td3tpcmLWMBP2FD0XBMWkaKrzzoatemrOiYs87N5F9Rlj7mI2NoQ3b2TuRZol8XHHKtvE3o
lCvLFtV8jQinOUq2S7mi57LKPfOTWpwEb5tNUk/UEltvMiNYygJEAFhQkiCgKtY+Begu/3eDULQN
HI4PC0jmDdEtydY7nMQ/bszmwshrnO+d4KL/weDjtPEzjRPSLFwqohE1PlMadZoKz6lDGlUqvlMy
zbOyYcn+mzAERB1HsieGQb/nXRUvX1lYx5eyoNssOYMWaUBGgc0ze622v3WHR1QEE1dpiouOevCS
I2sLEz843CHQ88hDN0uLmAJ9sYoN18wz94WJC0RMdED0pJBZmjG6Mr/+YgoI+ivl9mdjPQCV7+7i
KUOo/cTafFO1DN0U4G7AKIojGl5jmuw/7QyPJemeHjQkmyDdth8ipcMUtL7V9WjNvMgR2g9XFf5J
xrvnwE9ver2U5b1boFle1JyOJL9Y10Pxw0l4fjdpjSP2qe/oaGbfMj9MDDBovGUmOyf7d8kC8ot2
U9Rg/s3zu9/ItedrUNzXQzaCnUHMTdywmD/rrvO2MMQqECTZWSDLKt5PwUQvTPNSWm/pvnWyGuD8
hfXBzR6P7UV6OR8/hwml9mbq2zCmd/TohffdkJm1jCH9OgmQ2emm5ewz10izU5kkYv8om9iMsMpI
DD/CCZNdo5VQvnXQHERe42otokvmMPHc1c0+ibkWye1mtIdp317XQaFeoYOs335A/Oq+cMSR8ACt
PS6PvQG66qRUXl/H0K+yjmeo543MLrGechMlCRojo6IYpncA9UyQvUEe2ti9jyniOWwpWMChQa30
is4C1H1YwAhyshttqDQdpei+yJ3x7feIIE5KkfYUKlnJcoSWYfbV22Z/ALqfZx/1I0t3YAya68Vq
lkcFzPs8PcsbwXH6UOf5uNvf5DgV3Co2LCW58vzYCUTnFOf2YIR/FcJVcVAMMPMTDPcLCYaY06ze
S75CuJzTM42D7rqGHH8am2ByxdOZgJ9NwoAIiaRk5hecLVwlOFLmQLViFPi3m35DKNpA8XN9noxL
m276MFDU0RiKVe/PfUQAJllwFoXxukepH9Byvtkttyiq6XKJfo83BMjOlmIPfG2KaCs1z+9A0qGC
28gEeNDFeNGLSQsESjijGS/J1cKYDjr9hnY1b/bXPM28YKjR7H+Y2XNeU43GnZYWOXeNe6A3NlkK
/OHPeez+WPk4gNgnzNrGNLlYgBtn2xu0C6+9hEFqvQEArnP3BcVGgnOjDFiUVGJ90zICtbE9l6bC
OV8m2VJzU/McCcol0zxp7V5FEK5NPD7nXgwX9sSI4sMN/F9o1jzeasEkCvZffD2/1MQbcNPf/XhW
N6rbM7U4clc7JoslTIysJtiL4bkWKmOAS7y9Tr6ToA+JLtuwMLjwxTbDut2x3A6Q6d43JspT83O6
M8/R26a66pkrT1zypt6kJfvzv/EM0cWgWqCF3o+aU6IUUkKDDSDtsNMkEMwA+BxzQOKde1g4gYb4
juq6qFkAs9qRHP9Vhk2ZXqotu9Zn54jRiJHnOBcrNJkLGlug/pSe4uRQg7MSQbIPQv5pyQeE68cZ
qvJg7zMFcwrfHZt0ISf1M/pP1DijK72Ng8qnOVUMLnk8UUx6FzYIqLI2Uo/6XU0tEob5A1KNhobs
ZUxBhAfe630M19h4wfMWjX2+Yl95YQO2iUyIxF3vB4gO/ofdEIdMzi7+iqycTiWRQDJC1n42TjCl
wQvoLYKtnVNKnM7Ix/2xjacwnx6oA69Co8j8nV/Mx2ks+pKaXGdxyLKfeJ+mL9k4vcJlPHXaaL6G
GlZnKsH1vbQtXO0aQuD4TG5a0F0i/RuYKX6TpxFr5e46LwsnQUTPdbGByhKINCyUvWfXr8t3cpdB
pdUrpYvW9Og61bMrfeiRUZYPSQByfG7/xCB1R0XukND4/0kd4Sk6BHCc4CiScynMzFPKNkrEaQ6m
B4XPT3YwvnKOhuUILAN5fJ0PdA0qeuWFzmZODhJNtSinQ2yxCay5Z2mgaUa9vAfZ3+ziFFPGGJy5
h/C0x+NMt6zRmTVjNsek7Q0Dw2cJ5yJRnObqc9zky9R1l7pZgPImooXHBdhhWbUoUQ5/bVXprzYL
ukcf7kFWyqlGY6BHBvR6otVAI9ot8RUdXa2DeT+x9Ldc1gb9a8GZbU35pd0Mh1Pr6V2fmLfMiZA+
znjGG2d2rDCSZAdKeYK5bEV2xvyhiT6UEQy5C5QI+iheAavXhGGqyZwZ3RMizUHyYCcaHFrkhyUk
591YXQqVzkasixffPZZlLqRTArWtGy/8q0lREY1Yd7Ko2g3Sv+q3BJFa6sooSy800NpV5r6e43Y1
BlVK/LjbgX6SvzZvbVW0R2R8FQ0n6ArzRQ4RqJ5WXDL48lnncpiLGFYlVELPv22LzdDvhI47FknD
S0aPd7WmDxTc8n1elY7ONhKpKMX2zEJEYjCANjPeBv/akDkY8qwn1QVjwttGMYORbrh66eQdYSD1
AxDRmn7JnFPVNYvHK0S1D7AbjXOzrlBAXBBPgigUij+aoEXRi1yCGChLs20j6eFSF74EHuGfCirb
oY4t1iVXbOzB82wgGM4iUHshFnvI9XASBhQ1ISqWXpNNuz9sRPwsa5nMPwADa7CBQy+7N7lmBgs4
mBhhcIQRH+LydfBymHg98+jfCU9/FJHxe+jIMRZqvlo/M/s/zO9cHDGd6IGK35ahOIlIjJHoK/L3
UxMPTwz6eVQEBeT3eVtwpxGB2qqIlQn7zaMXlY2iOCkw7x7QhAOdzTgsbLIaHPmjJo5i35PEf8oX
hoZbunvI/ivGVMd/fvGNt+4U0WDof6E0H/KshU0lOyBR31VeWOi+HZOuTF1FJ060Hg4oxkDzguNw
F3F2cQgQFUu5bFzWI+iQzavrSSgu1E5fbYIz3ilize0b2+9O7r29ZOUof/pfayXum/DP8VAbrbHE
xxPW5W2HEciNZmSBJgekA5RgLM22PJLKX2p1BrVy0ss7UiPIr03M3hyCiy3YmT+mtHJQKG6uRlCi
X2jHsyRF/LnVz06lg1a/1KC6BeammHlJRrhs+NNGC2fvPsfJCJbRDlaYFC5b9z2ZYFDoxo5OzDru
IQZ3bpjh6oCNreKsLl6hJzqUt5hBe4B3WErEn23Z/dPX6KY7NBXSZGFX7N49cZKVhlO0xAsAcPFN
tfXk2P2+gokyEn8d4lyyU6ddyDqJHM3jiQA0bizLUKpmzyLMjHLrnVp4Tl/hmGYi3Ps09Nd1mRuT
mIAOKmj0sph/QXbCJApR6yKXSWA6GpoXRiDq1VDpo4sccxbfXVFLsBhPz4bolviyeDS0DAYLaWw4
n9RgWFvaAyCyXnVksR1mekC5oAMvzjp4OSobs+dSWCV9fv8fQzm0IaxccUvyq7clynAlI7ZjePNZ
hOfXC0SK+ruvQ2RtWvmM3jxMcpnT/HeEoKvqu4oXoC5N+yOGZGUEpZxjmuFSPAl+mIwPlCy8Gpwy
JBZjD1ywvRJw5pq+P5oYI7vDIDXwyKr/fRPGZt8Qermgry2WSjLnploSJeoRjPWkZfdP1Dj8iZWG
5OX+xKY8/s1gjebHzowDw9rs1DpwlG/J/LzAU+2AVBXCaiJWmtoK8NlW6CcEb6NnEAp6rWM4XX+j
wBKJlEvvwYskIl6Zt5wsydR5+aYlJdFfkgcJ477x3svsmoUwY0AxzdT1boR+pOa6lc+G0sm1lcVT
dfyU8LdoNb+9pfZna2+YnXOX7HjscFENrXs3/Nsw0knXJTDCpctWy0+BWIoe27k3bfa1d+Y0n8k2
CzyCozVtNCuFQcYcctXlKzMXydhS9gydhh/PxlnOqLGjXEvGJ5YYADS8XsRvYAkxrG8Bt4RflVqp
RuTNdOjLNUgFaTS2ERc8Qaz7WQkbyR5gqDcpmQAp/NY+h6smALlo+GnTfq4cwI7fyEKGJRazAsVF
IDsqLObvnXNJ5rXqkxj8RtpboAYHXl6x1kcEBmJ4FY1/D8evTYqyRqKSrO4ZY2yukAasMbJXAu5k
TaSGc5UDJ7C+6u6sXqBgSs5HdQmIdAu4zSl0oNKNXmVIAEEFuxJM1lkkuIG7+HT/oFVdYMFy42yV
oUOglSka6d8SvTtN0HOIsEAgpDxM8ftzNsoHzLJKGNUbUS22MV1E0/BtzJKPov3wZhIOZGsr2fff
LdcxpahtCEcwOIqOAqVGqq2yPkOYHsaU8C21Q9ipXrsrMuQzz1t7TE+OGbXuEm04tixxYAR18rub
GqOG/czcnGgznpL7pcjfic6Y5Fp2TWUbguM0dIppjmdYO0SoSjwFsk+VdZrsJQEuG3A+31gJ0iVE
RDmCNHf6zfFdBW+IpxydFifXq7+svPo0eWw0U/i9owP/9nl6R0Ca0/5wVtnEqyGrqkyqqVpkBodu
Hf1yTyirb0o+M1Wg5aN5+3zIT1GNPhSeRfFN6EDoui4ign3Co/qVXRw9T2keVSwsAigsfBfJJQPK
5GXePFrvOwD1qMKg3KjNNyJyyM4Q0DRr2WvHHhaujntc1GB+S76JoF5oN2F01Tr/qYVYfgE+uTiB
zbNCNCuze7zam3pwqsmHbnoytZYdu3OKCfzbHFsQq611K+SCsSeTuBSA7yr/jugr4bHnvbkbb3UJ
xgcxbzOIU7P9jGJ1U9c/EXidSgK8twnFNUsqWHRWm7wvW6SIePAia2nkg/sTs4JG2zV99j9RNDsq
jXnHl6BftFHwazTYRAWEoV64Lv0u7iBGrMjITsaTsFaysGN/sm9Q8MVp9OI9gkpcPbq8edtgbfDu
fgz9HPum/FnucIhcLN0kdLu4uXxZBpTuUa8CgQhgH6+/dRv28Nt/Det3pL81csZYLfFAcUDHyxch
WC9MfFAFHQGuhQGa3FnofcMFnwVFT9Yv09HCBN9jRKWq7xFPa1R3ry0NCSX8ESVGDyulvyi0YlFt
YcNCf4IUmsCHB6IkLw2zrcfcyFVazZn1v7pXl/qXYjr7IhNUVE5VHF8NBK/mEvMzIDz/2MSu2Qk0
8VVKQ2dX2usJIcsBYd8M61hA7aChNxRbg6kjngRotVufNlBUwYbBHuNQSt5BSOYU6LNyY3MtT+D/
Ql/cI0VmUq4B7vqC4Ts3R8qKMSKUfYD+1mUIVUxljV/YZHu8e6hVRmbXjPzujOhBADoRdl1C6hnu
gKNjWqvCDZEz7qnuYWv6/PBQ0WcW6T1xWVmCsiwgQXIFyNFg4JhZ5Fb/3N3YDjrmu6OWEwSufvvL
+4S6wYFv5DnsuCyHNswRGrRWX1giAztGfUplzlroPurf1E1sX7uMT7W9C+d8IkCBbzzarJhJmaGH
LzhUvVUgaKFIkva8zsXCx6N+dnkGTW1gM3gzrfm5AixKBqJMvPQRLiTCUN2aQlJzXruekM4lz9tf
PlumWJ1w0mhVEmTnTo4NQGr8iR4btYa0kOhFwTSLQMfXGfpHdd+DHyCXAIdCK7H3p2ywdcw1JC3I
6jw411osvvTQ7+ZDvDZtnPoXCcVWJZkylo3oOjWBzM+TvE5A3JYXNTM9NCO03+qkiZbHrcS9VyNK
UrCgijg9lBwADiiAdHkUuiLi2/aRVMRR3po/VkpL+fDgRYhMXi0vgy85qMFb0ZYN+OdjDM0aBjxV
N8M393MC8Hvv1P6UP271FLoEkeIivSDEyYJmnMZ5k0rmrTu0rhiaVAuFJKyZIKi+8vK6PiuI6cnE
+uBGQf/tTyRNqfiCbE9eIVo/c74aNimkeDT/ORSZhlaU39LSKrlh9mJ0dNVpnrVZft7Z7doZQQD5
EP/K8+vxgqrztzl/oqu0I9GC3dG4zfD1HCMckeGojwlUWxbrmaiSWoc6UgsTnM4k/CfR5QbDB1Gf
MJQtaL5HOa4uOQ/id8lM3swmFl+uki9p6hesVosodogEgtod05f83te0IdEZ9h+npgAbVh+3Kio7
JlbQEYTeh+01WHjfE9QaTIMoJ0wE/W7HRBt75ZRstq9KcdZW03qSiAjuwZCyJ8Dqcld5IU3NkPSV
jut+KxsbOKn5tkSQrsd8UEQoMySu9IvVassAU2T/XT9YuImJz5sSRb/5XGqP6jlJJxOdjgr1asoH
a8GozChFbKPbJsW0NQm+Vmjw/VP3TgPc+Z0CawwmisKfJpmuv8GwU9iGOgza7vqVwDmU64Yu6ko8
rMrSDmf/knCSZElAbtEsG5+v11Qw1LTnqH9g7vkXnpKMyMwdNzNW1zeAE1aC3TruxVkLxnjWGgw0
pkIv2PRW9AqzGf/T7Rc9kW7ZlFCKdvaNIDbwyOnDhdToAcxi5BI/CU9097LnTlSbLrnmgC5YomWr
/9h3Y4AStAdGM55JDShqnrlSwxMhaqUBQTHVM8C6yAnsvwCotMtedeEh5LTnzUYIOoUaDeOqbfmY
pRvMe2lR/x8wAprvILMtzI81cY2DLfvpJnlFuXWc23nFF2TAv1cZL2ZEOOkKGKG5B/GucqclnFLD
qNhfg0Az9e1JVd69SirbFWoWg7X4Ntsv/dMxN0NtRvXTpQ7peUmeGvTgz1XiDagjBcbnqb/TaeTT
GAgmEVNDcLvMnUDMGH5/z1T1luOhThFBmU0Tfma0zdE9qIKKA2CD8TjDaMeUhCV0+v398KE+UoKl
qTvekWb9yLvqDxtC7NzJCBx9LAatvUYR/2mqj6tgo0qJh3vlguS8S84g/UhwOqCW4Yuqq8UJ3WPc
6FGY1dSFRrjXsz7iJRLRvB4BS/8JAird03KzwiT7it9c1PW5vCchxGgNPNsxG0prwGNEy0SQ969m
G+zPYFqzYKanQO+HJIu1WQX/HlW4pkxmJpAHWTPuHd0JalUsnt5+ex2S4e9HIOhIjUmkV7OA0B+8
yr+wrJEs4kVoNP3pGrKu2L17XTlZH6NNRdR7wX4loBeX3JXI22O/4TGtbA0vXK13aoI868DYyKLL
wX5SkvI+TANK6r4BN4RJNen0agVUdambrF1PHu5eAp78bYMXKvOZGOYP5gxtdY1l5X8hZUBQsi7K
U59HQ5wHNgbvX8kzjnoBC3K1kMVEIwVXX8GOq0Ujn6P08XOCjLeIdc9XE1Al8PY06iPvcgZq6g7b
BeEtu1BaX1ULNkO7XgZ8Ib8U+ADNUgCY4bKmFvpM+2OH6qPl+h0sQMkuUdi0ec145BYszHrYvzh5
z6Om8bwrmz+eOrflGOnsuWwcy6/ymRzKQpawZJ/mhnIT+rr3BTtTYpFoDit1K2+Xrrhz7+Opcr8b
V34crPYXh0xBZsVha7JOLLBB6Yq+JXmWvIA9nZWmvtuWcyS36Xw2agmo06JSkAn7/d6UwHga30bL
smxPrnvqFPF02F86vVQ23f+e+rdU/PgNiywUrngZ+ECgY0TrtiHCo6lJxW50YDJ5BmSOLL0EVDWl
MDlalL1B7kLQPtMWiadVHMJ6IFENFvuib4Ntqr4zxnrZsFlVdUyDunfGZ/HspAxM3WTksvngmHzl
KR6t3qCHlo5yf7TUszQN3dTdUELFFNo34wZrROfmE699c5dfdMELWIBcThZ1REgGC+dfoYNwHA3J
8ai9xRc9d9fvelQPW8t+sg+fAi/t5RcZ+C3lT8ZKHZSf+figAxPqF1Hv0l8NdKeYbez8ZllRN7Yq
iT8E0K4YNVj1NlVoAswlN8aPwgvzIO+MWReebC47EWKlf3k0v0ZA/LujTBfuzXtJscIN6rxlYV5K
tSZdczl5Ek1t3VJ+WAcQShJ/GYnyIOxbuAXjLZm1gc59gwuL2xzsdZHHFnwUGcCGKAXE5y8IZWbu
rVJInwagxvg569lQ3A+34WkwX2uH91G9Q/7qdj5ly3rPEdjIPR/ku/CX+w/zonECgAHspFYJM9W+
mGEvpvnaFX5WwYwH3g8zlSeBoPHy5cgSjYywnSZMAQtp/0zuy/v28arvyQBNrjtP/91iChV4JH0m
cProRGd6IAcp0CyLTHCJQYxs+286SbGAn05qjtcNT0KZE42gZ3XWNuxbF17Gr86/xeeyxbVmePO8
0IqFMhTE+/UijiW2TDMcjMIKuTnga3XTOE9RsXqSEGzFoZiE2LxzU7upzDarbUscYXIy/PVvft1M
eNrLsu2NcjfpTe+tJHzH35qLBrf4RBS8HOCepvMC0aKb/huy/3v/blRdbwjImVzN2Glg+f5sLPvT
iu9CwImbiQYMg9memxCT2W9NHQLVYhAvZVQHVeMUFdOeyTTWhBTV4/CrQVBCKkHGVopKXwA3OqZv
5Yum+y5N8LjCdCzvyua6YKtivpc2bI9QBm/H8s1O0wyWIaW1iEAO8WAqMUfeCCK83Jz4wqFfq0sd
RYmXSBPiHcBnz00yDRUHLk1sNEtyo54lBkW6ckmwBHjh+pxjBu6n5NN0n+prtDhOtGXc4FArCzWW
OFwIuCFu6aTJSH384cRTSj0/H7yxs8+PVqpLOJCByPW+TOnHHxQx+Vz3r8Mvi5awho/JxIZ9ttnO
naGTgKdL30Mgrn4yU4gg5xVs0fyT2U3EumHRZ4ty/pXf31X+w85nt410JlqTaQdmdj07Boyoljn0
+Yai4X18/Aen5QI+vWYb9kpHshyoKyz+fwO77wbpMuSdmzyc2mJy5Pu0+sqr4aIfYiXKY2SRV8gs
SkNmr8dexadfBtAgnRu8/Zy2M5jXL74NOgr35ONeqgPZRYho31DWAzFLcyd9BP8JBwxUtDy+GR0I
Jt+dfIcmFL1admpuNhrDXATKwNa8CZl2DhRof3EojZc47RaKS1MZ5PPVUr7sUN9HY6gClG+m0Ug8
mu/Jny18b0UvWR95Pflo2WTaCMyMSvVjUwW3G1qH+a9YLYkQ2Z91MQFJLl9mbOZQqS5YA514kqhr
11RDDtCiaDE1dnH55vGLI6Dv7EQAnQMpcy/09lpwlauXysOgGWN2dt6LiTAH61o/MbSxNhqFclsA
pdza9C1G7D5pPzR0+HQuNz2KXizK2v1uvNwcN/V47e2gTWs9gH0Zd2yBT1lpKNBx9xoLhFW/+tb5
xTq2Nwh45/AqX9jVJhYChEwForzdEib4yfFFgd0ilnGZQikS2HLwx6JH6vYNUWggDhR0wau2YFma
tP+bNf1EL886Zr/OEyqkxTSvzU+RcVKArp7nVlA5JFDyOuF5EzfpJIzKktyw4ebXstS559XbE31N
xWfl++FEFOM/SWJCKulPtK0VmT4JDRXF4oiAQwocMWH4XDnbOCO+UQCHJNMrktB/qPyTq8duOlYI
FOM80cP4HA8L8kNRRmpjCiwpGREWGU205t76IkhvBjs6g7eDvoh2W5/QnWx7opKw0x7AJN2+C2g/
Ch+DbQPvRhELnmyJHTHmlxwa9Fw1QXNw6+UwGYCmaW+OTwFF5dgIfyNjqqz46ezevuxdSP1isaPr
OYt1Aj6QDWGZg8pRF8FhvAtOhNUm0Zrg8eM4yymQUmO3lCZ+ArFb0OPYxbX0YslcrxIuRR5EqnAK
iFKR+3yRFQLnCJF+YlfWaCxua2u7ODGuKPwmJiQTfGGbTbuac+TmpZmqMHfGkwmR+M8OKBytmDhD
K7gEkR66jqSgLiNRMLFSrl+0FTxjYG0H+IOKU5K2hYHIPuppoQxu/BM4eeSMNQc8T9kMtrd8cpxX
WIdDMC24/oYSRW/JnRmUc1VP/gbChgGQVP+uzp13Oo2N3cDQYJ+io8JPSX5aEMaib7b+uNHI9Vmi
PT6Sx2bS9KgMcbIx6rvp+HnhOvv01H+/59k0aorfemMsq/j5Jdn5XRIzSlLRgQtl3hlS3Qotx2XK
Wa3yXGYdBxbJp5mXuu6q19XG2a1pZxlsTGbiX82R3PoAcYO28bGnmJd96lMk93h+jTtRtBCBMiC9
s/mlQcV49PJLz+7kLFU5FXWq6Ua1JytgEwYuY21EF5Hskt8CNbu1AfeN4vR52AR1LWjYhs0huv4G
VSiJzHQFQ8MKSHrpqVmjY/bfMHTk6VNTrSXjoR28rkQtdd0mXwo8WhKocR/9Hz1R5m9x0nvgc3rG
mgYoIDiQRwr7ro+4iXDfGIvc2iq75GMYL9zDKKadB7piIHwo/Z0eaMMazg8K6gEdXC9htEBA5MSs
fAXUoynoMfoltLqK6UHiaO2Sk/0lvVTQJKiWlhfr5JneU+YmtYt9eu8FZHXTN2nWiubSAVPNgghw
J97aVp72LeL6A+6yYVWFn70k2e7IzQlvw84CO4dFUY5920PExSlJaWI14PsQc8WpjyLi4CySmBn2
wp/CcA/edzXUfcxSbyFuZ4YtajSMxNnro6Rqc44L9npA+qnnSfM+uKuX4QUYCl0zhc8rnZrHPFuj
uGZmMJF11xD9jz7sCjoPPxrFaZrSwNUCwGSBzY8Vw+5KyN9KrelUdbE0XjsWJehx7AX7H181W8aA
Adw9f/NP7eyF4uMJ6RthvzoYh0p4SoFhs/ZQ6vZ3BwF2PX3Xp7f2pB/rdGWfPRkaeF0PNzR4qqiy
TRKWVzwH3g0OocvD0GIPPASagejiIOlzjqhhHSPe5dy8hT/NWTutuVo8EJ5owfvcH7isp+RjQTAE
t1gjoGmdk3DRG63i1qUwjWvMHDy5sFzE2emOMawABFkMUq+9MOytFpAIc7GDVmR+66BLwH/R9oEx
ahYwa7f3cNG/l415vQf/zU0216ERW+BEHjbIietXBk4hWZED2paohKa4CFDX2oXSKoC9xoiFJ68D
1Q9uf+y4xyNrnjWHnhKoXYoSsdSLLjsk/glXF2CqC5KFInRV5vawFfAJMwjhM7xO2iMnGRQbiZd0
Vh8aZrhY3ExG+CTTlhMS4V9YiEGTOy3Q8S2i1gYEbaPNyo3ZTiYCbV/TLZo0LKQB+7v7hwa+WH1L
u3g8JtabJKtAizihlMiRo2sEZh+59rdUgpymPa8EbA6FUlBIfTh+0NNKOvLH/gZ/XfhxP37poHCU
z0kZSgArN67VQsqoDowqVNGr6D6ApY7E9JA1m2YF4BH09DIXRkWpCMKhqLgR0eRcfoGiG9/fbSrX
dQwK0f+yyY+3LyWoZkQukVpKB/9ao0PZlaV+6TTxN9xNWko2TiXcAZ1fCf1QVECBoL2ItyEoV51H
KLbTo8mhaeCCq9o74XUCYmLC0MYdXHAIBgj0T7a2SCEH0nGfHy2gt9FI2ytTMgQtjYXqnQzfhg73
7cQ0ghsEDqUyO/mCe8a6OFB8IgB1TuYsGqHlpnwivZAvYwSUGlopcMw83Rbq3V7xDvpIZDElMQ5+
vxqqGOAPIKSApmMMrffZRKSTRqyKrQ7Po398EPOi75qOBQLXkboYWBZ2S/I/MMGLlg41cnNc+Ykt
R9Hv8BE/HCsarBc7eI6u7/9Js5SOjvWLkF9HeqhvznF1Sg/GCCvoUQTrrSOpgmH6RN7DDD5QpuOr
P3PtmQmyLZfkYN2BNOG+BdE1YC1OhdGsLa0LceRTswPnpmWQw+dRA1hVSqY+5gc0bt0zHwYYpuyt
zg/Fn2f6XQGumUR5Fq9EfKtk1hhQM8K1rUnzWM3fiFffhnTenY3iTXhavnZkI/W13/KSlntiSXh3
gaUp3Fixns0RRlE2U7927bIVg/YqzuQT3FrPAjQRGPu/0Gw9aAcAxtch9n4l9v7KdMlvKxFeA3RU
jWyvnnj+bCLMfirk0n2v3TnOBhmQulRVTxfB6I8hHMdoiXkHNjwLWIzzur8Vn0tVWoC7MgrFiTeT
ZgnMgb9PLFJrUPpGdyYQ5WJrSIzymxK5MBM9qWz+2fMOoit0si72Z8275XU4Nnyf+5Hw1nkEbVDj
NgymRgAZny9xsCxuDyTA1x8317bc13h/skVjlmJLqQIs6q+5v7QmnbtyAZRgfAPuM3pLEPYh2x7i
n9NwCNK2FhgNgR1FW9tQ2URN9bEo7n8QsiOs65kClHkp2WctBaW1Cp6VFAXX1SvJShleLJTZfGnA
GWgQK5dL2DCu8wh/JAolsqMGL+6f+48x8MnN4nia4vQj0Gl6k6UEyS6aMsp2j+jwCmy1LMSFq5Od
9agSrWy/4QDVACoYAu0KW4H5ZmSJyOklMyZOXJThf2/Yv8YMXzSBchdnKqrXAoht7dfZXIhkLthR
iy5v/w5+++d2xKxdv24fUEpMdOATx+CM997wMCIa4xHo+jlFcgstDpYNIT9OkBOuNLi55MhceNnB
onspZ3LoRMWANjdoOgFJJMMmz39qcUw+1Oc4OPy1PXw7X0F8OK2MJVIgKRehMqGtTzgOxPRzgzF2
srcCh25w/ze/djOqypToBTF1L5VzaAHJNVRnaH0WZftSZIFQoE/zKGd/TAj3a6fpEGKT6rUYROYo
fH97B7lmzSTr8vrpyi+CRionIJVXmKK16HbBMwQXndNN7ApyreEM5mbc7P2zvr0OnGYdSWYSYPnW
sfUkXmghH5tCVqarDrrZTu7AMEDntL4kCsm4gTqdP15JJEP9DRsmE0hRTlnJj71WcJww39jtZwig
JxICyCwgTncIwCok6dHfVRRg8EM+GS2SlFxFTUb0cqKEkhHTg1VaRPlwJ+6UMaNQEjhsp13q1g/t
UsBLU7wuWI0H/7xr6Bfq0W5aZrYwbvHTH1rk6rPuHGginP/7D2DmJrK95RNmJQEoJOYfVC1oPmge
aEBKMlCdEcIwj2Y7yUvJS3ie2K7c+bIQiZrGwHQMQKDQWxoFyRU0squmWZxqx6k9CRWxv5OmKPeW
9l8HlWLq0cdmgf7ijdjSjblSd4tPfQvQBEWNSb5GbLZbFeAWovOFMc6qZDSNVBa3yAB7vur8ImXK
AGFOcHRTmwMGn3QAFePf4u7E0s1fyc7DvbgHK1ajD/0RHdoF7bsIKt8PzaXrBfZ1ujW5kJB32A9y
LBDp3CT5iV4roM0j+NXR+w8k1cMySXrthsCQW8oZ9GyabINc8nA8DFt35yCSZvH/T7A4bsFfx372
Q8YIKytwPir0Yoa7UschKTycN3iRWLWqtc7zF9rbR9EmS4/mGMmc7rnBJc4Nm90doB728A1LeMiy
AHGtOiJE8eKbLepHsFm2MUWrV/Ri7khBQ6bghXrsN0/9ng==
`pragma protect end_protected

