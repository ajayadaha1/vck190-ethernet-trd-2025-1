`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RrOblE+N+qIJxSW8DX3HlKoIR8i3b5/Q1epp13zuaL/Sr0ZUe6MdNQywZ/K2NfPkU8AGTkqYZaUI
BzXlCdodWSS8v86qM3cwZYTIymvLYQ+xXoTd0XWajVKsrXkIcwZs30ai7+P5OV+soZhqdnNjtGY0
2nxTfoyf63pZeMBtj+DWmydvc8e7dRVmQS9d/MzQUNPxz7f8ZVp7tYEz3VjaAKnyGx6sZpxN4QQY
RUP6FK/5IV2EK/p8KaQdBavkHOOQqIvZhAkLaxTSxcMd0DXNeQapvFJn3NvryueRBKFIZyL3NcIJ
1euH8bET136E9/mBk5y79Ne9/NZtQ8I/xnJI2A==
`pragma protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ZPm8TsbCbgY3d1ZBduuVPv19D1fXwy+2qDy+sTmiBypl7+TAUnjUF2d52uf+VwJPYbUYaQkd7bbL
tP0eqmb8pDdRwe5XS/a4b+CKfv2JwoaEBWt9BDWN9OMAGmdCNOAe43RGNujBIJ7+qSWRbjwrtIla
iRrBdVEe650sKT58YFWBDTyrNMW6TolSYZjAiCw3/B7hbfxr7ZzvyfKRLbI12KkBBivMjvVnd7+u
m6eZG+DpzkjutkOzGVRHx3X0ySy3Vu4bTB/AT3FutRmn/zkj0//pWUa4Ov8Zzxf2QPm5BNO4HIdY
eKmYfUbZ8e77OeMCrmjVMGjU2jzb+MG6ihF9wQ==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
VZ5pFILtbXU4Cp73V8lnfYwUyy1iCHqdcUHcmen134SQR24+DzvdK6mha7kaqbOZsboKe26swgZW
WqZN+MFq9w==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
lRY7rXGXeCruDlhvdxXdQ+BNwVLONYY0GAEN/9CkgDJFJWGNX59m327a3g0Q3VNCEvPV7cDY5mBB
iN2upmHUKXO3dyzS4wxCSFQyeDkSy4AAHnO5ebTjnPEAuhC6sN1Ypj+DJQXCk8cWPtN24++3AJOk
GM06El+GdMAsTMIX1y2CBNSngq/1NH5Spj9QjK/68OobafgaQz3WkdsroSq6ubqvfMz6yf9BnqTq
Zd6FCMlZF7eq4X9v9T4bOXJ96wyxNSMK4vZ/LjsVUydiHq2UZBNWHZkJPF6KOSjzi1pdIkZI/mTJ
cSCWzA0qcZIUZGmliAvqCd7eWdznvf5/tDcXRQ==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ANsd49vhYs2cfOxyRMxKyHxzi2VB+jCI0BWpGtUYhxtAIkzXAbCyCqPlEjoyAGa83sVBntmKbThR
ImF5R/X/c4NrpBunDYpjptXsnuMa1iaNafVaFlcN8a0BKK6nrdwjBfb13Xaxqric/8TRElmDEFGn
+3Qu5Sy3MSsF/1R0Em8=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kdimyzfoCuEFPizj5kpmwbCkoyvLzm+Zd7qZ2QFbflg41tODh66pkuGKYrTpxpQWuNRCoWNN1Mkh
0W9MI3tIQM2iQfmWM8V7WuoAr9Z9mdd0+OJW3/pRPCMEC03tntto1/wNBKRvM2iquO9xeIi1Rfzj
X3icEx1wXcVYU0H7yJbc4mWUlIDbXcPw2eCivcKWWjSePV5RDVlQ5G2kV3enhr3X8UpiefrGaGPF
p76FWVxsetxEu21obZvk/bB00yrvtqymPIkTn1Ca22ptTvqD9gcsOFDVKs8zaISzseHpbXnFVt3k
bsDq0QaYy4TzfTTdw+eRvL9MLhhXN8oEUNuJmA==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kx8QIu96mV5k9x0fZyNePjymbRR7xhfe0+IA8cvusZhORWS4VPtHvg0yt+xbA6JvRNTil3+1mdbc
UcBTqhTlzI+FZJjCH6YSUCuGJ9Iae2nWLnmwJ5dzdVSUZCfdWkufIKgWgCsvZUWrdmEcUEfny0rW
WC1qOvtE+OYddQ5OKA+nPODvPjxYFJWVYLQbEBcsNw899Cj5TU9SC6IsopcgeFCxXshcArWlnEmr
7mcIh+smFHorvqHHffJ1mrPtWuRSW8606YAlQpgqF4QQHDXwS9xJpMVPLn4+ha11ChkosAtWgpYC
QcJQwnDvjjo6Ejme2Fed2lcFjxOIpilVzik6RQ==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Gu/ChmsftRwJdFRsN6E6LaLXlBagxs9h/p4vkf34Y1jb7aQi5Ez3inMclpHVb24yhkqih6LqkEHO
nNjL848/Z5ZcFP/i78+FqDHT/vSWMDK6vaIGuXMJoDxcLHj6Y5p2Hdz/Age0GfmMbuBNiLvcf4My
b+V24ACbRbc2rZG68UI=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OCM3+2zE3VHEiOu9SHmcxLMwKvTRJ4WL3rpjCwAuzfxkA3i5vJqIUhXqADOsac09Y8mVBifLSd4O
9vmqhkcLJPBRoufM7+vvkwYo8fWvyfn6h21Ej1a5gfOLT/luI9U8qHWRofCCqR/mET2w1KUQr0rr
sEEtQuQjqD07Yy0e/z6L4msNOL94igOj1xiqqknfaVd8IzeCW1BBK2+8WbtlH4b3sMTfGv2RzV6V
htDXIMp/LnA8WGt3Jp+hn9uoMRgfgUI9tcb+m6wbqJ4Agr11VHzS3vK35hSJxVAHEFJEtpBOpZX1
H7tst+y0ggMCimFmor5UYpaX4pVXIa6SxAEn/w==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4544)
`pragma protect data_block
k34/+N0YVq+b3TeRsL8ghYNmg2GSn/7go8WkAvhuY+umenc7mDv0q9htzC+/0XT+EvWo/J4rjxG3
qSkEnYjT3c3/TbFz3GiVmcxhrB/ySqaaDqa29Kt2YIIrObQOXJw2EeeWe/2YW5LZ6KxizulwrC6/
L7NdjEIQG4dQwgopmXfVY56pqJHT61YSDFGPgbXy3srFTfcIxqaY7qWeUjP1ALvXjg/4tWvDE1XG
R2jKscKkdhLqUSyIRBMBAZjII3nQqUFWO2JuZl/9clzeq6gK9Ug7XKRyaC/w552hZ4ew9YQbxNIp
prrnuUUp8skLi+1uXc4sDGwHNYgxIzdIjlp6ln3OBpFsrQLQXhLbCRjlTQ85+gWjlV8BSTYlfNHu
xn+9En/nJ3UoAwJ4mpTv3jSIb4O5hTug01ANyYU49LiGbdyHmarN5POD+exvauSf/Y5OVMwi3HDM
S7K7WWQXzgWdqN5Q7AFj3oTc7ZczjQMLFV4dWgGSipT56Xo5aWaOLyYKh9YPDN8qwdprmcOKnMl0
rLwZAhZ3MLv7VEs3yaRvokUUE1fifq1zJewg/gvSMY1nqdqhg7Ag7RTTwAGTuDHZyXsOM9xqxS9f
NGuvQAXUOPM6WbQUqMFTGBg8wuv1FFYeyMNi4FnV0z0PdW75pH7Lknjdr1yEYFgz7fLLe4nSdtEq
RIo+5OhIAmOmWtlO2atXVw7TrwSnWpLNWa+NlXSeBjYH77r7pTlPxACnBeNe9UPx77exWJwE4Bg2
SxqtFplAAJngaB1ahUxDJPmgvBIYxlqTUorXjVwEQiHmfRsFv5JIm/56xfoPEk9ti94gNfv8UCvM
FqLttUTM6+bqeRUC9oFrBjPVbLAamLwKu9n6r2B7XCt6BPGlff8Xhk54PY8LkAFeB5KCIo++sI0C
VTdWtixPhwONY3GfYfuv+J+HyxDxlS1snESmvMFwG3/c5JXGtM1KuUGkYSmTvkdATgbsp4k0QZ6N
ZUn+WQ7rce570BLjrqRShFDynlWcdGuy3s8uPzyMpw6Zr4JQr+M4I5A5Fk3pGLOcOtcBb06inn0D
WvLCB4dH1Z7lSZZpbMUuHr6N61RJriI5FOaafSUoOXp//XcOSvFPJZrFk1ak7tI8cOgPewpO/poS
flVlAFATyMi0SEeV/gwsPDzdlp81Ey5KldUzVQ387iQEYbf8OYtNRGLDkqz/8GAbbi08R2AvQ+dG
Y3VqE4ONumE4D0Dy5p7K5A0yAOfLnmEpn3ocyoxaGbU2IoL8n35naWFMeWV72GKfALXW/OnyMx+P
JDdHQD38D7Iq6qG44xnUKsmzUv7qRew5HaaP8eZ2Vt4PyfHnxFZ01MxogsPIN3LwL1iUPsna5efN
TWsWO2WwEp5a+sZU6jXAuAEkwmDzMlBaJErwk8X5ASffLl+dYnnoXvRuoSZPkd8cyA3NX9d03S3x
3vBgVChBIY0Dq5VSDqwHCA5HBehMYCEAa4dEmLbDGt6JTQcd7tRkrKBEivY/+2NQGB/847mQXy1Z
fGXU5gstNRFCVD2Gaa0uBmWwJF5rEc9Q0hFsOkwNRtJ/dvkQlaRoHlaakqrknq9E+BfMDo89Goza
NVdhDtj+Y8CR8TwOgRsdRm7YbW2hd1nYCgKgMjg6tZ4WOimdGSQSTZm2f2qSU2m+8emfz4QkiiMo
xf4he9r2uC8FUUS7s020K9ikuiIZKgb7O0kKf+BrFMyU4SxAqA20wLD82RF8ywjVE7/bIfUAu5Iz
/3RX01vFxBO9qC+yNj36GVv3huAx+DP7f4IY9gL0De3EqH689lRo9QNUHIRKjqlC+NAs9GijaNv3
bMZ8eHEl/8pBrkgKxhgRZDOKL/lA6AAYkAB/HTP6Cm2mKHWhhZMfphlLq9ziaTaeyoqcWX7mw6NF
Rhp6k3vSKnsHNNP+G3sgVjFVb4JrrcAyVEOj5irW6Jr+qIYNuNylMck1ZwIoHevHfCAcHsqA6Oxb
brHwWyfI7diKBpI6Ewan4rnw6t7P9jFBFsD2e2WoUf/LotG4t0RaCEgDK1WO9UqxrUkSYgZsWQdV
peUrOmBw7h7dRCCmIp08h8Cnnv5jFqGoiq5X1pBJsSmkYohgnLP+ELqBDIAHQpnOfXqLJeB6JasQ
90cA0npRvqtB+yUozxhFY9kJ9aLjZNjl+zPfIhFqg1d6ORZqKPseT4OhO+fXqRsc1CLWXA15oBml
1uBAxq8UQuXacaJQiz/tyQRyCA3Wjrfahf+xF9vIDkhmVc0JsunYiHd0+PI8/bIHgyzqL/v/Mgzh
uCvLQulpg9PCPuwD4Nk9V/D3CqOqCMsrYm7YdwiWjboo43K/bht5BNJLoj8L2AHHa69Kb/luwFD+
szLHhWrn8SMfWiXsBxR+MKNAmWdIQziMFC5E3M2YGS6wbxFqoTJD7O6pPI7sbWU7QvV4V3QBPcvn
bfdGvwtnbIYIGV4AomYMlyiZnWBlCRRTkZOx3eIg5EmziZJpHkgMYSi3l+ooi9HfkQIROnhg/hDF
fkN5PAThbPiU7teU+/BakJqPpfhQStbyFEJnS7pegiYpgrpUNG04PJd/mRhPW1MM1bYFbsrcNbZJ
Jvj3kmGkDMzKTuOEUDL0aKr37kzEwTZ38l5/ogCEijplaI73FxvRxjw4y60AJjnRKO46QEl9TkPY
OLf84LOe5hi3zwE/6+NvqAARcwgDpbj76f3V+ysXlM526YxMFIYZXENewx00q/57waS+vcKZelLE
afhFJecKka71ZfDxXHmoQDJjEuaLRjHQMvtJFo4PK0rWpxDWyvLdd1gvfeVXvtD6xgg85j734VRX
RQ4bOetMe/kMJQG9YUwnp3etMGh6BhaHJJpukvKlsHVKdyUO6L6WlKLRLqdMC+YsA+9nz+Jw/eC4
Zo04TxlUpygUzu0ksAArAlZRnagUycIh3kQ5tJfGEMOja0MFZD8rJEX1scXIE9WvIFUK5qM0andn
ouTA4RTOmBStil319ewTbn24GY04cbQ0EoOd5x6c8aJMWr2AdjN2RfVOLlDGLy55tklBIIoDBSeB
l2RqmVUZxcJzPjC8pGkvNKshtTAIUT42YLNpIBT1fz7lpKRMJ/gH9JH+sct1Fz1rFxsaCkLihQNx
tEmaqrAF0INov3I14UmcAS3AXbU6rABltecABSRttXMS3KI/9fi8kOVkNseH1+hL1c+wksOL5yHO
ApiZbVb7nw4nEz/QnZ/xWfRLAzQ47tzh0aL6gscsJYO3IkYyva2dyA0JTF1DT24WrFuAVJlNwJVY
1kkK6Tvyk/zH8fnJ7rRcTjhU7PWPcy4uOZFsKl178dk2EGN2MQb51KGK9dv/lC6EvGZh4T5mvhk9
/hULFW3uU7akzn66ovwhvpcOov8eL1EpJnu0qQNhHHnZDgkwaiRLHS4aUzFdOPAdmzx9iU50qU7Y
avL9EA4ds55fxF6YLhE+8NoO/peH51fwbTOqVjpGaTw2jmRCSuZupY+diHDJHLZR0QmH2WdgcKn+
XXoIgIHfUeLtIBxQyiii75xvhBJY/1QQhNg5wSArIbtUv97oslIoGpCBN1ly1XyLJzDCjRQk/7kM
GC1LYST+hW1v9Jf/3cYaXy5M54iurh97pFk4PzgsxoNc2J5VC8vb3N36nYp4gLTxWBafrniT5ego
vUPWysLriEyMQ0+VGNoajfVPYPWCHpfMER8nU8Aj0jipz7yvUFckaTM4i2PPdFY4hNsmHd2wEGP8
Zi2eZjxzFm46lRZawBWfR2km2vFHvzrSuABhAdF9ryGNJfd1KjM+dsk6nYFfeFQG8wjU4gufHnex
dxqL68mmjDRCp1Y2pQ4kJPiTcTzn/51inGvm7Cc3oE8f8GvGOPz8f+/lVzNYB/pEyUfQ0LqiXB66
CghcZOzFLG6DkZYaSwWg1fyNVZ+1SR8KgWkDpd6B7c77O/xyoc7s5/FJDDZyqwR1QRR9xGcuf9TB
8d4wzRJ7H+J0WlubcDSk1EI9wVm0LuDKI0OmkBMNRGlNWMQxkdc8kiF3ZiyPmU09zg2CKRqGtqIz
owx0BWFitKtNnb8McQVkMsGZ+v7BgTqPDqP2rtVgAuSphM0jZPbiwUxfqSHq1kl1rhYhDSgFKsxv
L9CyQpXqE8q8zF6h5QtudCVLS/RvBhmPG8bouUTyF0QOphsRyvfHXzB/ZjOnUgFjVRgDEwwpWlnV
ZLCDdkyYekXGY7v1tk/xXAD3wxVIph/VPx6s5PtDpsfnXD/J5GtO9x/MwUShlkLS9Nx9sOHrcAcJ
k2L6KwLe2EDduu6hbF2A9Eblf3fAD4VtUKIio9kInZOL16iMx9LqVLhO1VdZqO3/R9THDpk+sUkW
BHRa5vlkxBjz4NlEcjSdY9sFxc3KXFN+z9uAzpOcFf0Ty+mvi0lL7K6f0WcsN/KfBhUkrY2zwrRs
N7eOz010+IMz3CaOjb+e9ZjPlo2pKyLG7r+cD44ke0TwH9Xr3TEuoHmNVykvnjqrwoHt1/dy69t1
maDoVE1e3d5y6aXQBzy2CEigR/c/eZTROvzo9O0dG+/3CnHjkah8AvrWGSbNAfOwZ3+woG1yFOW9
OOra8JyqtphyYjFv8u1Ut6sdr6NMMkPll2+zEg7FyPRmCxS3sZlAy34YvCoS7A276PlReQqwTPs5
7Pi6VcKVyGNTCD696VzK1etBXxdvbikIru3dDHSWgB27WS76L5j95sRSxsIECm0vfWiIEZPiuuUH
AlfauyFqPa06vKUEmyku69yzK6E5fYcSP8B9HS6tbMsUGe2hUS+XaUWl9wyv57EfBu1UNnYpt6lj
BkSKfeLZoEOQ7KVW802d5YiLu+amEmJD3Cyd9Uyjd5iszR1xXJJqcj6vCGqbG2gog/8QaiCRCqIY
Rz7b4YZDJ6qweVNEkOewQwTN1eclZ7Ix1axv/PepBOVY11iPZjK//9cKdVLFTHS6L6aJoLwGSraI
JZd76+74jSIWNwBS8vuApyiaki/uhWC0Ovlh33ml8AQdzAV/q3d+sFs8uClyOkWdkfOdCQEkcYmJ
DaP89Kql2EjeN/aEyUaWOR5LNGZbcsYrW/XEJDoQAvGVeBDsBLq35Y4q0GupFhJOv4MAP27F4BM6
is1nAV8vZi/iBRuY4WoRpe0aS9aRKTsE6cnS9GYdNqJft7JTwfSBup6rVgovYMygFsZc5407Gf6V
gVClHAe1mbDaarP+GhBMoZD2xS6qiPGyCjmOrubhqAIOhnL9sTrM0as3shGsFikSTYD96EPUmo+i
jstreK376aYfuedTOu0DFpS0N2KLJzzCnCxcLZCB9RsKCTb23/bXq30pBIL5tUGSKlOzk5RdGf6K
XfJp1llRAT7C4RplXNbzruOshIf7lYtMtU5MvMkGfAPoGTrp84n/fm7cigIGAySsYmP3tLpC67XO
+b+1FWnC+nxGDlOpqQWyoi3+ZMiXofzDxU6SicP/4t3QCDcjQb5AXZOwPNXfW4QuR8VB3i08Gx7c
SWUCWL0Hf22uaCvMlJbu5r3bN6/vbL4gFJGE2D2hhQLdOjiAostiN9/YCAzniHFGyHle8Qap9+bf
5hUbwhEpkFnmg1s0LyrrAAQT9SWSn/G5ZAd/FCKn7g/apGdVDgDIWASJr/YNaBmayMaJf9UMkoUU
YrbfhQM5lako/oZdvOSZOtDPWinbCvYVpNloFqe+3cP6jnT/3VKpgbmvMeiEZ4E0udMOnqIHiBby
k4yL10lBRGWbkMEnyanfRzww0d334xOfi4XckST9U1gjpRVemlr2Sce1nP79PmnadzeOPIBI1jaw
TQT8g4QYqnCUn1SehfkbjfIMYgbgpbkcQQjM6MyqluR83m0apOgxQU5zwRTSCFy54EIuaG7l5kqG
EkgbJOdKd4R5D7MD6o0/qVh54/zqQcsgWrCie4XEdeaqpzTIzcszh97HSlcOfnO2NUA9d3XnNxpk
gvdZIWukxVDXUHXiAeloVRhPkMRaRomFhwWlDJjFjE15d1kMIHobEz/tMKmwhk20aeitbis70qop
JvLDwxpQaFSKWjcERkwEODt7OeM2YPtqcT0JVlZsTxXRi/H8m7mf3Go=
`pragma protect end_protected

